magic
tech scmos
magscale 1 2
timestamp 1744796300
<< metal1 >>
rect 824 2006 830 2014
rect 838 2006 844 2014
rect 852 2006 858 2014
rect 866 2006 872 2014
rect 204 1937 227 1943
rect 164 1897 179 1903
rect 493 1897 540 1903
rect 573 1903 579 1923
rect 573 1897 611 1903
rect 1149 1897 1171 1903
rect 1188 1897 1203 1903
rect 29 1877 51 1883
rect 148 1877 163 1883
rect 516 1877 531 1883
rect 2445 1877 2460 1883
rect 724 1857 755 1863
rect 1124 1856 1132 1864
rect 2004 1857 2019 1863
rect 2580 1857 2595 1863
rect 2426 1836 2428 1844
rect 2520 1836 2524 1844
rect 2072 1806 2078 1814
rect 2086 1806 2092 1814
rect 2100 1806 2106 1814
rect 2114 1806 2120 1814
rect 538 1776 540 1784
rect 125 1757 147 1763
rect 573 1743 579 1763
rect 701 1757 716 1763
rect 564 1737 579 1743
rect 733 1737 748 1743
rect 1684 1737 1699 1743
rect 1796 1737 1811 1743
rect 2084 1737 2179 1743
rect 77 1717 115 1723
rect 132 1717 163 1723
rect 221 1717 252 1723
rect 420 1717 451 1723
rect 605 1717 620 1723
rect 637 1717 675 1723
rect 797 1717 883 1723
rect 893 1717 931 1723
rect 925 1697 931 1717
rect 1662 1717 1676 1723
rect 1725 1717 1740 1723
rect 1997 1723 2003 1736
rect 1980 1717 2003 1723
rect 2061 1717 2188 1723
rect 1836 1712 1844 1716
rect 1980 1712 1988 1717
rect 2317 1723 2323 1743
rect 2317 1717 2376 1723
rect 2452 1717 2467 1723
rect 1773 1697 1795 1703
rect 2557 1697 2595 1703
rect 1844 1677 1875 1683
rect 2525 1677 2540 1683
rect 282 1636 284 1644
rect 410 1636 412 1644
rect 490 1636 492 1644
rect 596 1636 598 1644
rect 824 1606 830 1614
rect 838 1606 844 1614
rect 852 1606 858 1614
rect 866 1606 872 1614
rect 1252 1576 1254 1584
rect 1780 1536 1782 1544
rect 2516 1537 2540 1543
rect 29 1517 44 1523
rect 212 1497 227 1503
rect 477 1497 515 1503
rect 669 1497 691 1503
rect 797 1497 899 1503
rect 1277 1503 1283 1523
rect 1277 1497 1315 1503
rect 1748 1497 1772 1503
rect 1900 1503 1908 1508
rect 1892 1497 1908 1503
rect 2540 1503 2548 1508
rect 2540 1497 2578 1503
rect 148 1477 163 1483
rect 909 1477 963 1483
rect 1021 1477 1059 1483
rect 1332 1477 1363 1483
rect 1853 1477 1875 1483
rect 516 1457 531 1463
rect 580 1457 604 1463
rect 644 1457 659 1463
rect 1725 1457 1740 1463
rect 2052 1457 2099 1463
rect 890 1436 892 1444
rect 2509 1437 2524 1443
rect 2072 1406 2078 1414
rect 2086 1406 2092 1414
rect 2100 1406 2106 1414
rect 2114 1406 2120 1414
rect 1764 1376 1766 1384
rect 1005 1357 1020 1363
rect 1101 1344 1107 1363
rect 1716 1356 1724 1364
rect 61 1323 67 1343
rect 500 1337 531 1343
rect 989 1337 1020 1343
rect 1108 1337 1123 1343
rect 1709 1337 1747 1343
rect 52 1317 67 1323
rect 1156 1317 1171 1323
rect 1261 1317 1276 1323
rect 2061 1323 2067 1343
rect 2084 1337 2131 1343
rect 2141 1337 2156 1343
rect 2061 1317 2163 1323
rect 2237 1317 2275 1323
rect 1876 1297 1891 1303
rect 2269 1297 2275 1317
rect 2548 1317 2563 1323
rect 2308 1297 2323 1303
rect 909 1277 956 1283
rect 1869 1277 1908 1283
rect 1869 1257 1875 1277
rect 1172 1236 1174 1244
rect 2170 1236 2172 1244
rect 824 1206 830 1214
rect 838 1206 844 1214
rect 852 1206 858 1214
rect 866 1206 872 1214
rect 2148 1137 2163 1143
rect 2516 1137 2547 1143
rect 749 1097 787 1103
rect 925 1103 931 1123
rect 1044 1116 1052 1124
rect 1220 1116 1228 1124
rect 820 1097 883 1103
rect 893 1097 931 1103
rect 964 1097 979 1103
rect 1076 1097 1091 1103
rect 1268 1097 1283 1103
rect 1469 1097 1484 1103
rect 2365 1097 2396 1103
rect 708 1077 739 1083
rect 957 1077 995 1083
rect 1165 1077 1180 1083
rect 1309 1077 1324 1083
rect 1485 1077 1507 1083
rect 1485 1064 1491 1077
rect 2397 1077 2419 1083
rect 1341 1057 1356 1063
rect 2168 1036 2172 1044
rect 2072 1006 2078 1014
rect 2086 1006 2092 1014
rect 2100 1006 2106 1014
rect 2114 1006 2120 1014
rect 2141 977 2156 983
rect 356 937 387 943
rect 461 937 499 943
rect 1053 937 1068 943
rect 1101 943 1107 963
rect 1812 957 1827 963
rect 1101 937 1116 943
rect 1124 937 1139 943
rect 1837 937 1859 943
rect 1933 937 1964 943
rect 2237 937 2259 943
rect 397 917 435 923
rect 1060 917 1075 923
rect 1805 917 1820 923
rect 2013 917 2028 923
rect 2196 917 2211 923
rect 925 897 1004 903
rect 1028 896 1036 904
rect 1924 897 1939 903
rect 1988 898 1992 906
rect 1676 892 1684 896
rect 1677 877 1731 883
rect 1556 836 1558 844
rect 824 806 830 814
rect 838 806 844 814
rect 852 806 858 814
rect 866 806 872 814
rect 1002 736 1004 744
rect 2164 736 2166 744
rect 1860 716 1868 724
rect 397 697 435 703
rect 884 697 963 703
rect 1213 697 1228 703
rect 1309 697 1324 703
rect 1357 697 1395 703
rect 1924 697 1939 703
rect 2100 697 2163 703
rect 2413 697 2428 703
rect 2493 697 2515 703
rect 356 677 387 683
rect 1261 677 1299 683
rect 1805 677 1820 683
rect 2077 677 2140 683
rect 916 657 947 663
rect 1396 657 1411 663
rect 2077 657 2083 677
rect 2221 677 2259 683
rect 2324 677 2339 683
rect 2509 677 2515 697
rect 2589 677 2626 683
rect 1981 637 1996 643
rect 2072 606 2078 614
rect 2086 606 2092 614
rect 2100 606 2106 614
rect 2114 606 2120 614
rect 490 576 492 584
rect 1444 557 1459 563
rect 356 537 387 543
rect 509 537 547 543
rect 836 537 866 543
rect 1213 537 1251 543
rect 1316 537 1331 543
rect 1796 537 1811 543
rect 2388 537 2428 543
rect 2861 537 2876 543
rect 2700 524 2708 528
rect 397 517 435 523
rect 516 517 531 523
rect 605 517 636 523
rect 2125 517 2179 523
rect 2372 517 2396 523
rect 2404 517 2444 523
rect 2541 517 2556 523
rect 2868 517 2883 523
rect 2036 497 2076 503
rect 2317 497 2339 503
rect 2013 477 2100 483
rect 2013 457 2019 477
rect 2122 436 2124 444
rect 2925 437 2940 443
rect 824 406 830 414
rect 838 406 844 414
rect 852 406 858 414
rect 866 406 872 414
rect 397 297 435 303
rect 1060 297 1091 303
rect 2221 297 2275 303
rect 2308 297 2323 303
rect 2461 297 2515 303
rect 356 277 387 283
rect 964 277 1043 283
rect 1213 277 1228 283
rect 2164 277 2211 283
rect 2349 277 2364 283
rect 2072 206 2078 214
rect 2086 206 2092 214
rect 2100 206 2106 214
rect 2114 206 2120 214
rect 2660 176 2662 184
rect 404 157 419 163
rect 1373 157 1388 163
rect 356 137 387 143
rect 452 137 467 143
rect 1060 137 1091 143
rect 1357 137 1388 143
rect 452 117 467 123
rect 461 97 467 117
rect 1261 117 1276 123
rect 1309 117 1347 123
rect 824 6 830 14
rect 838 6 844 14
rect 852 6 858 14
rect 866 6 872 14
<< m2contact >>
rect 830 2006 838 2014
rect 844 2006 852 2014
rect 858 2006 866 2014
rect 396 1976 404 1984
rect 668 1976 676 1984
rect 1036 1976 1044 1984
rect 1228 1976 1236 1984
rect 1548 1976 1556 1984
rect 1628 1976 1636 1984
rect 2268 1958 2276 1966
rect 2844 1958 2852 1966
rect 28 1936 36 1944
rect 140 1936 148 1944
rect 300 1936 308 1944
rect 332 1936 340 1944
rect 92 1916 100 1924
rect 204 1916 212 1924
rect 268 1916 276 1924
rect 316 1916 324 1924
rect 412 1916 420 1924
rect 460 1916 468 1924
rect 60 1896 68 1904
rect 140 1896 148 1904
rect 156 1896 164 1904
rect 220 1896 228 1904
rect 284 1896 292 1904
rect 364 1896 372 1904
rect 540 1896 548 1904
rect 588 1916 596 1924
rect 1036 1916 1044 1924
rect 1548 1916 1556 1924
rect 1628 1916 1636 1924
rect 2268 1912 2276 1920
rect 2348 1916 2356 1924
rect 2412 1916 2420 1924
rect 2844 1912 2852 1920
rect 636 1896 644 1904
rect 1036 1896 1044 1904
rect 1084 1896 1092 1904
rect 1180 1896 1188 1904
rect 1258 1896 1266 1904
rect 1340 1896 1348 1904
rect 1644 1896 1652 1904
rect 1836 1896 1844 1904
rect 2092 1896 2100 1904
rect 2284 1896 2292 1904
rect 2860 1896 2868 1904
rect 140 1876 148 1884
rect 444 1876 452 1884
rect 476 1876 484 1884
rect 508 1876 516 1884
rect 620 1876 628 1884
rect 940 1876 948 1884
rect 1100 1876 1108 1884
rect 1132 1876 1140 1884
rect 1452 1876 1460 1884
rect 1724 1876 1732 1884
rect 2204 1876 2212 1884
rect 2380 1876 2388 1884
rect 2460 1876 2468 1884
rect 2556 1876 2564 1884
rect 2780 1876 2788 1884
rect 12 1856 20 1864
rect 108 1856 116 1864
rect 252 1856 260 1864
rect 348 1856 356 1864
rect 428 1856 436 1864
rect 716 1856 724 1864
rect 908 1856 916 1864
rect 1132 1856 1140 1864
rect 1180 1856 1188 1864
rect 1420 1856 1428 1864
rect 1756 1856 1764 1864
rect 1996 1856 2004 1864
rect 2172 1856 2180 1864
rect 2396 1856 2404 1864
rect 2572 1856 2580 1864
rect 2748 1856 2756 1864
rect 92 1836 100 1844
rect 204 1836 212 1844
rect 572 1836 580 1844
rect 1916 1836 1924 1844
rect 2428 1836 2436 1844
rect 2524 1836 2532 1844
rect 2078 1806 2086 1814
rect 2092 1806 2100 1814
rect 2106 1806 2114 1814
rect 44 1776 52 1784
rect 540 1776 548 1784
rect 684 1776 692 1784
rect 2028 1776 2036 1784
rect 2172 1776 2180 1784
rect 2268 1776 2276 1784
rect 2492 1776 2500 1784
rect 2588 1776 2596 1784
rect 12 1756 20 1764
rect 460 1756 468 1764
rect 508 1756 516 1764
rect 92 1736 100 1744
rect 188 1736 196 1744
rect 204 1736 212 1744
rect 300 1736 308 1744
rect 332 1736 340 1744
rect 364 1736 372 1744
rect 428 1736 436 1744
rect 556 1736 564 1744
rect 716 1756 724 1764
rect 748 1756 756 1764
rect 1164 1756 1172 1764
rect 1500 1756 1508 1764
rect 1756 1756 1764 1764
rect 1900 1756 1908 1764
rect 1916 1756 1924 1764
rect 2156 1756 2164 1764
rect 2748 1756 2756 1764
rect 620 1736 628 1744
rect 748 1736 756 1744
rect 764 1736 772 1744
rect 860 1736 868 1744
rect 940 1736 948 1744
rect 972 1736 980 1744
rect 1196 1736 1204 1744
rect 1468 1736 1476 1744
rect 1676 1736 1684 1744
rect 1740 1736 1748 1744
rect 1788 1736 1796 1744
rect 1820 1736 1828 1744
rect 1948 1736 1956 1744
rect 1996 1736 2004 1744
rect 2012 1736 2020 1744
rect 2076 1736 2084 1744
rect 124 1716 132 1724
rect 172 1716 180 1724
rect 252 1716 260 1724
rect 284 1716 292 1724
rect 348 1716 356 1724
rect 412 1716 420 1724
rect 476 1716 484 1724
rect 620 1716 628 1724
rect 28 1696 36 1704
rect 44 1696 52 1704
rect 140 1696 148 1704
rect 236 1696 244 1704
rect 252 1696 260 1704
rect 316 1696 324 1704
rect 380 1696 388 1704
rect 524 1696 532 1704
rect 652 1696 660 1704
rect 908 1696 916 1704
rect 956 1716 964 1724
rect 1292 1716 1300 1724
rect 1372 1716 1380 1724
rect 1676 1716 1684 1724
rect 1740 1716 1748 1724
rect 1836 1716 1844 1724
rect 1852 1716 1860 1724
rect 1964 1716 1972 1724
rect 2188 1716 2196 1724
rect 2300 1716 2308 1724
rect 2332 1736 2340 1744
rect 2428 1736 2436 1744
rect 2444 1736 2452 1744
rect 2780 1736 2788 1744
rect 2444 1716 2452 1724
rect 2540 1716 2548 1724
rect 2860 1716 2868 1724
rect 1260 1700 1268 1708
rect 1404 1700 1412 1708
rect 1692 1696 1700 1704
rect 2028 1696 2036 1704
rect 2268 1696 2276 1704
rect 2492 1696 2500 1704
rect 2844 1700 2852 1708
rect 1836 1676 1844 1684
rect 1948 1676 1956 1684
rect 2540 1676 2548 1684
rect 1404 1654 1412 1662
rect 1852 1656 1860 1664
rect 2844 1654 2852 1662
rect 284 1636 292 1644
rect 412 1636 420 1644
rect 492 1636 500 1644
rect 588 1636 596 1644
rect 1004 1636 1012 1644
rect 1260 1636 1268 1644
rect 1772 1636 1780 1644
rect 2508 1636 2516 1644
rect 2588 1636 2596 1644
rect 830 1606 838 1614
rect 844 1606 852 1614
rect 858 1606 866 1614
rect 60 1576 68 1584
rect 268 1576 276 1584
rect 604 1576 612 1584
rect 1148 1576 1156 1584
rect 1244 1576 1252 1584
rect 1436 1576 1444 1584
rect 1916 1576 1924 1584
rect 2428 1576 2436 1584
rect 2572 1576 2580 1584
rect 2348 1558 2356 1566
rect 2828 1558 2836 1566
rect 316 1536 324 1544
rect 1164 1536 1172 1544
rect 1196 1536 1204 1544
rect 1772 1536 1780 1544
rect 1932 1536 1940 1544
rect 2444 1536 2452 1544
rect 2508 1536 2516 1544
rect 2540 1536 2548 1544
rect 44 1516 52 1524
rect 76 1516 84 1524
rect 92 1516 100 1524
rect 204 1516 212 1524
rect 428 1516 436 1524
rect 492 1516 500 1524
rect 588 1516 596 1524
rect 764 1516 772 1524
rect 876 1516 884 1524
rect 988 1516 996 1524
rect 1132 1516 1140 1524
rect 108 1496 116 1504
rect 124 1496 132 1504
rect 172 1496 180 1504
rect 204 1496 212 1504
rect 316 1496 324 1504
rect 332 1496 340 1504
rect 460 1496 468 1504
rect 604 1496 612 1504
rect 748 1496 756 1504
rect 780 1496 788 1504
rect 1036 1496 1044 1504
rect 1068 1496 1076 1504
rect 1100 1496 1108 1504
rect 1148 1496 1156 1504
rect 1244 1496 1252 1504
rect 1292 1516 1300 1524
rect 1436 1516 1444 1524
rect 1804 1516 1812 1524
rect 1820 1516 1828 1524
rect 1996 1516 2004 1524
rect 2348 1512 2356 1520
rect 2476 1516 2484 1524
rect 2828 1512 2836 1520
rect 1388 1496 1396 1504
rect 1436 1496 1444 1504
rect 1740 1496 1748 1504
rect 1772 1496 1780 1504
rect 1884 1496 1892 1504
rect 1916 1496 1924 1504
rect 1964 1496 1972 1504
rect 2284 1496 2292 1504
rect 2396 1496 2404 1504
rect 2460 1496 2468 1504
rect 2524 1496 2532 1504
rect 2652 1496 2660 1504
rect 2860 1496 2868 1504
rect 44 1476 52 1484
rect 140 1476 148 1484
rect 252 1476 260 1484
rect 348 1476 356 1484
rect 396 1476 404 1484
rect 444 1476 452 1484
rect 556 1476 564 1484
rect 700 1476 708 1484
rect 732 1476 740 1484
rect 812 1476 820 1484
rect 1084 1476 1092 1484
rect 1116 1476 1124 1484
rect 1212 1476 1220 1484
rect 1228 1476 1236 1484
rect 1324 1476 1332 1484
rect 1532 1476 1540 1484
rect 1756 1476 1764 1484
rect 2284 1476 2292 1484
rect 2764 1476 2772 1484
rect 12 1456 20 1464
rect 236 1456 244 1464
rect 284 1456 292 1464
rect 380 1456 388 1464
rect 508 1456 516 1464
rect 540 1456 548 1464
rect 604 1456 612 1464
rect 636 1456 644 1464
rect 924 1456 932 1464
rect 1004 1456 1012 1464
rect 1564 1456 1572 1464
rect 1740 1456 1748 1464
rect 1884 1456 1892 1464
rect 2044 1456 2052 1464
rect 2252 1456 2260 1464
rect 2732 1456 2740 1464
rect 204 1436 212 1444
rect 364 1436 372 1444
rect 428 1436 436 1444
rect 716 1436 724 1444
rect 892 1436 900 1444
rect 988 1436 996 1444
rect 1820 1436 1828 1444
rect 2524 1436 2532 1444
rect 2572 1436 2580 1444
rect 2078 1406 2086 1414
rect 2092 1406 2100 1414
rect 2106 1406 2114 1414
rect 76 1376 84 1384
rect 476 1376 484 1384
rect 1036 1376 1044 1384
rect 1084 1376 1092 1384
rect 1660 1376 1668 1384
rect 1756 1376 1764 1384
rect 1900 1376 1908 1384
rect 2588 1376 2596 1384
rect 268 1356 276 1364
rect 492 1356 500 1364
rect 748 1356 756 1364
rect 1020 1356 1028 1364
rect 1452 1356 1460 1364
rect 1724 1356 1732 1364
rect 2188 1356 2196 1364
rect 2284 1356 2292 1364
rect 2332 1356 2340 1364
rect 2780 1356 2788 1364
rect 44 1316 52 1324
rect 300 1336 308 1344
rect 460 1336 468 1344
rect 492 1336 500 1344
rect 556 1336 564 1344
rect 716 1336 724 1344
rect 1020 1336 1028 1344
rect 1100 1336 1108 1344
rect 1148 1336 1156 1344
rect 1228 1336 1236 1344
rect 1484 1336 1492 1344
rect 1692 1336 1700 1344
rect 1948 1336 1956 1344
rect 106 1316 114 1324
rect 380 1316 388 1324
rect 444 1316 452 1324
rect 508 1316 516 1324
rect 572 1316 580 1324
rect 828 1316 836 1324
rect 1052 1316 1060 1324
rect 1068 1316 1076 1324
rect 1148 1316 1156 1324
rect 1276 1316 1284 1324
rect 1372 1316 1380 1324
rect 1628 1316 1636 1324
rect 1788 1316 1796 1324
rect 1868 1316 1876 1324
rect 1932 1316 1940 1324
rect 2028 1316 2036 1324
rect 2076 1336 2084 1344
rect 2156 1336 2164 1344
rect 2204 1336 2212 1344
rect 2300 1336 2308 1344
rect 2412 1336 2420 1344
rect 2460 1336 2468 1344
rect 2540 1336 2548 1344
rect 2812 1336 2820 1344
rect 2220 1316 2228 1324
rect 396 1296 404 1304
rect 652 1300 660 1308
rect 1132 1296 1140 1304
rect 1196 1296 1204 1304
rect 1548 1300 1556 1308
rect 1724 1296 1732 1304
rect 1772 1296 1780 1304
rect 1868 1296 1876 1304
rect 2252 1296 2260 1304
rect 2348 1316 2356 1324
rect 2428 1316 2436 1324
rect 2492 1316 2500 1324
rect 2540 1316 2548 1324
rect 2700 1316 2708 1324
rect 2300 1296 2308 1304
rect 2460 1296 2468 1304
rect 2476 1296 2484 1304
rect 2588 1296 2596 1304
rect 2620 1296 2628 1304
rect 2876 1300 2884 1308
rect 12 1276 20 1284
rect 956 1276 964 1284
rect 1820 1276 1828 1284
rect 1852 1276 1860 1284
rect 652 1254 660 1262
rect 1548 1254 1556 1262
rect 2380 1276 2388 1284
rect 2508 1276 2516 1284
rect 2492 1256 2500 1264
rect 396 1236 404 1244
rect 556 1236 564 1244
rect 1164 1236 1172 1244
rect 1292 1236 1300 1244
rect 2172 1236 2180 1244
rect 2876 1236 2884 1244
rect 830 1206 838 1214
rect 844 1206 852 1214
rect 858 1206 866 1214
rect 44 1176 52 1184
rect 332 1176 340 1184
rect 396 1176 404 1184
rect 1084 1176 1092 1184
rect 1516 1176 1524 1184
rect 1596 1176 1604 1184
rect 1772 1176 1780 1184
rect 1916 1176 1924 1184
rect 1980 1176 1988 1184
rect 2844 1158 2852 1166
rect 684 1136 692 1144
rect 2140 1136 2148 1144
rect 2508 1136 2516 1144
rect 44 1116 52 1124
rect 396 1116 404 1124
rect 764 1116 772 1124
rect 252 1096 260 1104
rect 380 1096 388 1104
rect 604 1096 612 1104
rect 796 1096 804 1104
rect 812 1096 820 1104
rect 1020 1116 1028 1124
rect 1052 1116 1060 1124
rect 1196 1116 1204 1124
rect 1228 1116 1236 1124
rect 1308 1116 1316 1124
rect 2124 1116 2132 1124
rect 2492 1116 2500 1124
rect 2508 1116 2516 1124
rect 2556 1116 2564 1124
rect 2844 1112 2852 1120
rect 956 1096 964 1104
rect 1052 1096 1060 1104
rect 1068 1096 1076 1104
rect 1132 1096 1140 1104
rect 1228 1096 1236 1104
rect 1260 1096 1268 1104
rect 1356 1096 1364 1104
rect 1388 1096 1396 1104
rect 1420 1096 1428 1104
rect 1452 1096 1460 1104
rect 1484 1096 1492 1104
rect 1948 1096 1956 1104
rect 2012 1096 2020 1104
rect 2140 1096 2148 1104
rect 2188 1096 2196 1104
rect 2236 1096 2244 1104
rect 2396 1096 2404 1104
rect 2460 1096 2468 1104
rect 2524 1096 2532 1104
rect 2586 1096 2594 1104
rect 2668 1096 2676 1104
rect 2876 1096 2884 1104
rect 140 1076 148 1084
rect 492 1076 500 1084
rect 700 1076 708 1084
rect 812 1076 820 1084
rect 1068 1076 1076 1084
rect 1180 1076 1188 1084
rect 1244 1076 1252 1084
rect 1260 1076 1268 1084
rect 1324 1076 1332 1084
rect 1372 1076 1380 1084
rect 1404 1076 1412 1084
rect 1436 1076 1444 1084
rect 1708 1076 1716 1084
rect 1724 1076 1732 1084
rect 1756 1076 1764 1084
rect 1804 1076 1812 1084
rect 2300 1076 2308 1084
rect 2428 1076 2436 1084
rect 2444 1076 2452 1084
rect 2492 1076 2500 1084
rect 2780 1076 2788 1084
rect 172 1056 180 1064
rect 524 1056 532 1064
rect 716 1056 724 1064
rect 908 1056 916 1064
rect 1004 1056 1012 1064
rect 1116 1056 1124 1064
rect 1324 1056 1332 1064
rect 1356 1056 1364 1064
rect 1484 1056 1492 1064
rect 2220 1056 2228 1064
rect 2268 1056 2276 1064
rect 2748 1056 2756 1064
rect 924 1036 932 1044
rect 1980 1036 1988 1044
rect 2044 1036 2052 1044
rect 2172 1036 2180 1044
rect 2204 1036 2212 1044
rect 2412 1036 2420 1044
rect 2078 1006 2086 1014
rect 2092 1006 2100 1014
rect 2106 1006 2114 1014
rect 492 976 500 984
rect 1196 976 1204 984
rect 1596 976 1604 984
rect 2156 976 2164 984
rect 172 956 180 964
rect 364 956 372 964
rect 556 956 564 964
rect 764 956 772 964
rect 140 936 148 944
rect 348 936 356 944
rect 732 936 740 944
rect 1068 936 1076 944
rect 1084 936 1092 944
rect 1356 956 1364 964
rect 1772 956 1780 964
rect 1804 956 1812 964
rect 1916 956 1924 964
rect 2044 956 2052 964
rect 2316 956 2324 964
rect 2764 956 2772 964
rect 1116 936 1124 944
rect 1388 936 1396 944
rect 1532 936 1540 944
rect 1644 936 1652 944
rect 1788 936 1796 944
rect 1884 936 1892 944
rect 1964 936 1972 944
rect 2028 936 2036 944
rect 2188 936 2196 944
rect 2476 936 2484 944
rect 2508 936 2516 944
rect 2796 936 2804 944
rect 252 916 260 924
rect 444 916 452 924
rect 524 916 532 924
rect 588 916 596 924
rect 620 916 628 924
rect 844 916 852 924
rect 1036 916 1044 924
rect 1052 916 1060 924
rect 1164 916 1172 924
rect 1484 916 1492 924
rect 1548 916 1556 924
rect 1628 916 1636 924
rect 1692 916 1700 924
rect 1756 916 1764 924
rect 1820 916 1828 924
rect 1868 916 1876 924
rect 2028 916 2036 924
rect 2156 916 2164 924
rect 2188 916 2196 924
rect 2268 916 2276 924
rect 2332 916 2340 924
rect 2428 916 2436 924
rect 2492 916 2500 924
rect 2540 916 2548 924
rect 2876 916 2884 924
rect 44 896 52 904
rect 412 896 420 904
rect 668 900 676 908
rect 1004 896 1012 904
rect 1036 896 1044 904
rect 1452 900 1460 908
rect 1580 896 1588 904
rect 1596 896 1604 904
rect 1676 896 1684 904
rect 1708 896 1716 904
rect 1900 896 1908 904
rect 1916 896 1924 904
rect 1980 898 1988 906
rect 2172 896 2180 904
rect 2236 896 2244 904
rect 2284 896 2292 904
rect 2300 896 2308 904
rect 2444 896 2452 904
rect 2460 896 2468 904
rect 2524 896 2532 904
rect 2604 896 2612 904
rect 2860 900 2868 908
rect 1660 876 1668 884
rect 2140 876 2148 884
rect 2364 876 2372 884
rect 2412 876 2420 884
rect 2556 876 2564 884
rect 332 856 340 864
rect 1452 854 1460 862
rect 2428 856 2436 864
rect 2860 854 2868 862
rect 44 836 52 844
rect 668 836 676 844
rect 1548 836 1556 844
rect 1724 836 1732 844
rect 2540 836 2548 844
rect 830 806 838 814
rect 844 806 852 814
rect 858 806 866 814
rect 44 776 52 784
rect 572 776 580 784
rect 1180 776 1188 784
rect 1452 776 1460 784
rect 1804 776 1812 784
rect 1900 776 1908 784
rect 2620 776 2628 784
rect 2908 776 2916 784
rect 1708 758 1716 766
rect 332 736 340 744
rect 1004 736 1012 744
rect 1980 736 1988 744
rect 2156 736 2164 744
rect 2188 736 2196 744
rect 44 716 52 724
rect 412 716 420 724
rect 572 716 580 724
rect 1036 716 1044 724
rect 1228 716 1236 724
rect 1372 716 1380 724
rect 1708 712 1716 720
rect 1820 716 1828 724
rect 1852 716 1860 724
rect 1884 716 1892 724
rect 2012 716 2020 724
rect 2428 716 2436 724
rect 2556 716 2564 724
rect 2908 716 2916 724
rect 252 696 260 704
rect 444 696 452 704
rect 476 696 484 704
rect 604 696 612 704
rect 876 696 884 704
rect 972 696 980 704
rect 988 696 996 704
rect 1068 696 1076 704
rect 1100 696 1108 704
rect 1228 696 1236 704
rect 1324 696 1332 704
rect 1340 696 1348 704
rect 1532 696 1540 704
rect 1740 696 1748 704
rect 1852 696 1860 704
rect 1916 696 1924 704
rect 1996 696 2004 704
rect 2028 696 2036 704
rect 2092 696 2100 704
rect 2204 696 2212 704
rect 2268 696 2276 704
rect 2300 696 2308 704
rect 2316 696 2324 704
rect 2396 696 2404 704
rect 2428 696 2436 704
rect 2460 696 2468 704
rect 140 676 148 684
rect 348 676 356 684
rect 460 676 468 684
rect 508 676 516 684
rect 668 676 676 684
rect 862 676 870 684
rect 1036 676 1044 684
rect 1084 676 1092 684
rect 1132 676 1140 684
rect 1324 676 1332 684
rect 1644 676 1652 684
rect 1788 676 1796 684
rect 1820 676 1828 684
rect 1836 676 1844 684
rect 1916 676 1924 684
rect 2044 676 2052 684
rect 172 656 180 664
rect 364 656 372 664
rect 700 656 708 664
rect 908 656 916 664
rect 1020 656 1028 664
rect 1276 656 1284 664
rect 1388 656 1396 664
rect 1420 656 1428 664
rect 1612 656 1620 664
rect 1948 656 1956 664
rect 2140 676 2148 684
rect 2316 676 2324 684
rect 2380 676 2388 684
rect 2444 676 2452 684
rect 2524 696 2532 704
rect 2876 696 2884 704
rect 2556 676 2564 684
rect 2812 676 2820 684
rect 2236 656 2244 664
rect 2348 656 2356 664
rect 2364 656 2372 664
rect 2780 656 2788 664
rect 1228 636 1236 644
rect 1452 636 1460 644
rect 1900 636 1908 644
rect 1996 636 2004 644
rect 2060 636 2068 644
rect 2572 636 2580 644
rect 2078 606 2086 614
rect 2092 606 2100 614
rect 2106 606 2114 614
rect 492 576 500 584
rect 1292 576 1300 584
rect 1404 576 1412 584
rect 2828 576 2836 584
rect 172 556 180 564
rect 364 556 372 564
rect 556 556 564 564
rect 716 556 724 564
rect 732 556 740 564
rect 748 556 756 564
rect 1020 556 1028 564
rect 1228 556 1236 564
rect 1436 556 1444 564
rect 1612 556 1620 564
rect 2252 556 2260 564
rect 2284 556 2292 564
rect 2300 556 2308 564
rect 2332 556 2340 564
rect 2412 556 2420 564
rect 2556 556 2564 564
rect 2924 556 2932 564
rect 140 536 148 544
rect 348 536 356 544
rect 460 536 468 544
rect 572 536 580 544
rect 828 536 836 544
rect 1052 536 1060 544
rect 1308 536 1316 544
rect 1644 536 1652 544
rect 1788 536 1796 544
rect 1964 536 1972 544
rect 2140 536 2148 544
rect 2188 536 2196 544
rect 2236 536 2244 544
rect 2316 536 2324 544
rect 2380 536 2388 544
rect 2428 536 2436 544
rect 2876 536 2884 544
rect 2892 536 2900 544
rect 252 516 260 524
rect 444 516 452 524
rect 508 516 516 524
rect 588 516 596 524
rect 636 516 644 524
rect 684 516 692 524
rect 700 516 708 524
rect 764 516 772 524
rect 780 516 788 524
rect 940 516 948 524
rect 1148 516 1156 524
rect 1196 516 1204 524
rect 1260 516 1268 524
rect 1356 516 1364 524
rect 1372 516 1380 524
rect 1740 516 1748 524
rect 1836 516 1844 524
rect 1884 516 1892 524
rect 1932 516 1940 524
rect 1948 516 1956 524
rect 2012 516 2020 524
rect 2364 516 2372 524
rect 2396 516 2404 524
rect 2444 516 2452 524
rect 2524 516 2532 524
rect 2556 516 2564 524
rect 2588 516 2596 524
rect 2652 516 2660 524
rect 2700 516 2708 524
rect 2716 516 2724 524
rect 2748 516 2756 524
rect 2780 516 2788 524
rect 2860 516 2868 524
rect 44 496 52 504
rect 412 496 420 504
rect 476 496 484 504
rect 620 496 628 504
rect 652 496 660 504
rect 1148 496 1156 504
rect 1708 500 1716 508
rect 1900 496 1908 504
rect 1916 496 1924 504
rect 2028 496 2036 504
rect 2076 496 2084 504
rect 2156 496 2164 504
rect 2572 496 2580 504
rect 2636 496 2644 504
rect 2764 496 2772 504
rect 2828 496 2836 504
rect 1868 476 1876 484
rect 1996 476 2004 484
rect 332 456 340 464
rect 1708 454 1716 462
rect 1884 456 1892 464
rect 2604 476 2612 484
rect 2668 476 2676 484
rect 2796 476 2804 484
rect 2268 456 2276 464
rect 44 436 52 444
rect 1148 436 1156 444
rect 1404 436 1412 444
rect 2124 436 2132 444
rect 2204 436 2212 444
rect 2492 436 2500 444
rect 2588 436 2596 444
rect 2652 436 2660 444
rect 2780 436 2788 444
rect 2940 436 2948 444
rect 830 406 838 414
rect 844 406 852 414
rect 858 406 866 414
rect 44 376 52 384
rect 492 376 500 384
rect 652 376 660 384
rect 1196 376 1204 384
rect 1244 376 1252 384
rect 1420 376 1428 384
rect 1772 376 1780 384
rect 1836 376 1844 384
rect 2124 376 2132 384
rect 2636 376 2644 384
rect 2924 376 2932 384
rect 1516 358 1524 366
rect 2428 356 2436 364
rect 332 336 340 344
rect 940 336 948 344
rect 1164 336 1172 344
rect 2412 336 2420 344
rect 44 316 52 324
rect 412 316 420 324
rect 652 316 660 324
rect 1068 316 1076 324
rect 1180 316 1188 324
rect 1516 312 1524 320
rect 1836 316 1844 324
rect 2236 316 2244 324
rect 2300 316 2308 324
rect 2380 316 2388 324
rect 2476 316 2484 324
rect 2540 316 2548 324
rect 2636 316 2644 324
rect 252 296 260 304
rect 444 296 452 304
rect 636 296 644 304
rect 860 296 868 304
rect 1020 296 1028 304
rect 1052 296 1060 304
rect 1100 296 1108 304
rect 1164 296 1172 304
rect 1692 296 1700 304
rect 1852 296 1860 304
rect 2300 296 2308 304
rect 2364 296 2372 304
rect 2396 296 2404 304
rect 2556 296 2564 304
rect 2572 296 2580 304
rect 2636 296 2644 304
rect 2844 296 2852 304
rect 140 276 148 284
rect 348 276 356 284
rect 460 276 468 284
rect 604 276 612 284
rect 748 276 756 284
rect 956 276 964 284
rect 1116 276 1124 284
rect 1228 276 1236 284
rect 1292 276 1300 284
rect 1308 276 1316 284
rect 1580 276 1588 284
rect 1932 276 1940 284
rect 2156 276 2164 284
rect 2252 276 2260 284
rect 2284 276 2292 284
rect 2364 276 2372 284
rect 2444 276 2452 284
rect 2492 276 2500 284
rect 2732 276 2740 284
rect 172 256 180 264
rect 364 256 372 264
rect 780 256 788 264
rect 1052 256 1060 264
rect 1132 256 1140 264
rect 1612 256 1620 264
rect 1964 256 1972 264
rect 2316 256 2324 264
rect 2588 256 2596 264
rect 2764 256 2772 264
rect 2540 236 2548 244
rect 2078 206 2086 214
rect 2092 206 2100 214
rect 2106 206 2114 214
rect 428 176 436 184
rect 540 176 548 184
rect 1244 176 1252 184
rect 1852 176 1860 184
rect 2204 176 2212 184
rect 2300 176 2308 184
rect 2652 176 2660 184
rect 2684 176 2692 184
rect 2860 176 2868 184
rect 172 156 180 164
rect 364 156 372 164
rect 396 156 404 164
rect 876 156 884 164
rect 1068 156 1076 164
rect 1228 156 1236 164
rect 1388 156 1396 164
rect 1564 156 1572 164
rect 2044 156 2052 164
rect 2460 156 2468 164
rect 140 136 148 144
rect 348 136 356 144
rect 444 136 452 144
rect 508 136 516 144
rect 652 136 660 144
rect 844 136 852 144
rect 1052 136 1060 144
rect 1164 136 1172 144
rect 1276 136 1284 144
rect 1388 136 1396 144
rect 1596 136 1604 144
rect 1740 136 1748 144
rect 2012 136 2020 144
rect 2492 136 2500 144
rect 2636 136 2644 144
rect 2732 136 2740 144
rect 2812 136 2820 144
rect 252 116 260 124
rect 334 116 342 124
rect 396 116 404 124
rect 444 116 452 124
rect 44 96 52 104
rect 492 116 500 124
rect 956 116 964 124
rect 1100 116 1108 124
rect 1148 116 1156 124
rect 1180 116 1188 124
rect 1196 116 1204 124
rect 1276 116 1284 124
rect 1292 116 1300 124
rect 1692 116 1700 124
rect 2124 116 2132 124
rect 2380 116 2388 124
rect 2588 116 2596 124
rect 2716 116 2724 124
rect 2764 116 2772 124
rect 2828 116 2836 124
rect 2892 116 2900 124
rect 780 100 788 108
rect 1036 96 1044 104
rect 1212 96 1220 104
rect 1324 96 1332 104
rect 1404 96 1412 104
rect 1660 100 1668 108
rect 1916 96 1924 104
rect 2556 100 2564 108
rect 2668 96 2676 104
rect 2684 96 2692 104
rect 2748 96 2756 104
rect 2860 96 2868 104
rect 2876 96 2884 104
rect 2780 76 2788 84
rect 2908 76 2916 84
rect 1660 54 1668 62
rect 2764 56 2772 64
rect 2892 56 2900 64
rect 44 36 52 44
rect 780 36 788 44
rect 1116 36 1124 44
rect 1916 36 1924 44
rect 2556 36 2564 44
rect 830 6 838 14
rect 844 6 852 14
rect 858 6 866 14
<< metal2 >>
rect 381 2037 403 2043
rect 493 2037 515 2043
rect 605 2037 627 2043
rect 653 2037 675 2043
rect 781 2037 787 2043
rect 397 1984 403 2037
rect 13 1864 19 1936
rect 141 1923 147 1936
rect 141 1917 163 1923
rect 157 1904 163 1917
rect 61 1884 67 1896
rect 93 1764 99 1836
rect 13 1704 19 1756
rect 45 1704 51 1756
rect 61 1584 67 1736
rect 157 1724 163 1896
rect 221 1884 227 1896
rect 269 1864 275 1916
rect 285 1904 291 1936
rect 189 1764 195 1856
rect 205 1804 211 1836
rect 189 1744 195 1756
rect 301 1744 307 1756
rect 173 1724 179 1736
rect 77 1524 83 1676
rect 109 1504 115 1556
rect 125 1504 131 1716
rect 205 1704 211 1736
rect 237 1704 243 1716
rect 285 1703 291 1716
rect 317 1704 323 1796
rect 333 1744 339 1756
rect 365 1724 371 1736
rect 381 1704 387 1916
rect 413 1843 419 1916
rect 445 1884 451 1896
rect 509 1884 515 2037
rect 413 1837 435 1843
rect 429 1744 435 1837
rect 477 1804 483 1876
rect 541 1784 547 1896
rect 269 1697 291 1703
rect 269 1664 275 1697
rect 269 1584 275 1656
rect 285 1504 291 1636
rect 333 1504 339 1576
rect 141 1484 147 1496
rect 45 1324 51 1476
rect 237 1464 243 1496
rect 285 1464 291 1476
rect 317 1464 323 1496
rect 349 1484 355 1496
rect 397 1484 403 1736
rect 429 1704 435 1736
rect 461 1684 467 1756
rect 477 1724 483 1756
rect 557 1744 563 1896
rect 621 1884 627 2037
rect 669 1984 675 2037
rect 1085 2023 1091 2043
rect 1149 2037 1155 2043
rect 1245 2037 1251 2043
rect 1069 2017 1091 2023
rect 824 2006 830 2014
rect 838 2006 844 2014
rect 852 2006 858 2014
rect 866 2006 872 2014
rect 1037 1924 1043 1976
rect 573 1764 579 1836
rect 685 1784 691 1916
rect 717 1864 723 1896
rect 717 1764 723 1856
rect 909 1824 915 1856
rect 749 1764 755 1776
rect 765 1744 771 1796
rect 941 1744 947 1876
rect 621 1724 627 1736
rect 861 1724 867 1736
rect 1037 1724 1043 1896
rect 413 1584 419 1636
rect 429 1524 435 1536
rect 493 1524 499 1636
rect 525 1544 531 1696
rect 589 1644 595 1676
rect 589 1524 595 1636
rect 605 1584 611 1716
rect 621 1664 627 1716
rect 957 1704 963 1716
rect 445 1484 451 1516
rect 461 1464 467 1496
rect 541 1464 547 1516
rect 605 1504 611 1556
rect 77 1384 83 1456
rect 317 1404 323 1456
rect 13 1284 19 1296
rect 45 1124 51 1176
rect 141 1084 147 1196
rect 173 1064 179 1356
rect 301 1344 307 1376
rect 365 1364 371 1436
rect 381 1344 387 1456
rect 381 1104 387 1316
rect 397 1244 403 1296
rect 397 1124 403 1176
rect 173 964 179 1056
rect 45 844 51 896
rect 45 724 51 776
rect 173 664 179 956
rect 253 924 259 1096
rect 253 704 259 916
rect 413 864 419 896
rect 429 884 435 1436
rect 445 1324 451 1396
rect 509 1363 515 1456
rect 557 1404 563 1476
rect 500 1357 515 1363
rect 557 1344 563 1356
rect 573 1324 579 1356
rect 621 1324 627 1656
rect 653 1404 659 1696
rect 824 1606 830 1614
rect 838 1606 844 1614
rect 852 1606 858 1614
rect 866 1606 872 1614
rect 733 1484 739 1536
rect 877 1524 883 1536
rect 765 1504 771 1516
rect 781 1504 787 1516
rect 749 1484 755 1496
rect 925 1484 931 1516
rect 957 1504 963 1696
rect 1005 1583 1011 1636
rect 1005 1577 1027 1583
rect 701 1444 707 1476
rect 813 1464 819 1476
rect 925 1464 931 1476
rect 989 1463 995 1516
rect 989 1457 1004 1463
rect 717 1364 723 1436
rect 653 1262 659 1300
rect 717 1284 723 1336
rect 557 1204 563 1236
rect 824 1206 830 1214
rect 838 1206 844 1214
rect 852 1206 858 1214
rect 866 1206 872 1214
rect 685 1124 691 1136
rect 813 1104 819 1116
rect 612 1097 627 1103
rect 525 1044 531 1056
rect 493 984 499 1016
rect 557 964 563 996
rect 333 724 339 736
rect 445 704 451 916
rect 525 884 531 916
rect 477 704 483 876
rect 589 784 595 916
rect 573 724 579 776
rect 365 564 371 656
rect 45 444 51 496
rect 45 324 51 376
rect 173 264 179 556
rect 253 304 259 516
rect 365 504 371 556
rect 445 524 451 696
rect 461 544 467 676
rect 509 563 515 656
rect 493 557 515 563
rect 333 324 339 336
rect 173 244 179 256
rect 173 164 179 236
rect 253 124 259 296
rect 365 264 371 496
rect 413 463 419 496
rect 404 457 419 463
rect 365 164 371 256
rect 397 164 403 456
rect 429 184 435 476
rect 445 304 451 516
rect 445 164 451 296
rect 461 284 467 536
rect 477 484 483 496
rect 493 384 499 557
rect 557 544 563 556
rect 573 544 579 676
rect 589 564 595 776
rect 605 704 611 1096
rect 621 924 627 1097
rect 717 1004 723 1056
rect 765 964 771 1036
rect 813 1024 819 1076
rect 909 1064 915 1136
rect 957 1124 963 1276
rect 957 1104 963 1116
rect 989 1104 995 1436
rect 1021 1364 1027 1577
rect 1069 1524 1075 2017
rect 1277 2004 1283 2043
rect 1485 2037 1491 2043
rect 1549 2037 1555 2043
rect 2221 2037 2227 2043
rect 2525 2037 2531 2043
rect 1229 1984 1235 1996
rect 1549 1924 1555 1976
rect 1629 1924 1635 1976
rect 2269 1920 2275 1958
rect 1085 1704 1091 1896
rect 1101 1884 1107 1916
rect 2845 1920 2851 1958
rect 1181 1864 1187 1896
rect 1165 1764 1171 1816
rect 1149 1584 1155 1636
rect 1197 1624 1203 1736
rect 1341 1724 1347 1896
rect 1453 1864 1459 1876
rect 1421 1824 1427 1856
rect 1501 1764 1507 1816
rect 1261 1644 1267 1700
rect 1245 1584 1251 1616
rect 1101 1504 1107 1536
rect 1037 1384 1043 1496
rect 1069 1444 1075 1496
rect 1117 1464 1123 1476
rect 1085 1384 1091 1456
rect 1117 1344 1123 1456
rect 1133 1343 1139 1516
rect 1245 1504 1251 1516
rect 1293 1484 1299 1516
rect 1373 1504 1379 1716
rect 1405 1662 1411 1700
rect 1501 1624 1507 1756
rect 1645 1743 1651 1896
rect 1645 1737 1667 1743
rect 1437 1524 1443 1576
rect 1325 1484 1331 1496
rect 1133 1337 1148 1343
rect 1069 1324 1075 1336
rect 1053 1304 1059 1316
rect 1085 1184 1091 1276
rect 1060 1117 1075 1123
rect 1069 1104 1075 1117
rect 669 844 675 900
rect 765 824 771 956
rect 845 904 851 916
rect 669 684 675 696
rect 701 664 707 816
rect 824 806 830 814
rect 838 806 844 814
rect 852 806 858 814
rect 866 806 872 814
rect 749 564 755 576
rect 509 324 515 516
rect 621 504 627 536
rect 685 524 691 556
rect 733 504 739 556
rect 781 524 787 576
rect 909 504 915 656
rect 925 584 931 1036
rect 1005 904 1011 1056
rect 1037 924 1043 1096
rect 1069 1064 1075 1076
rect 1069 1024 1075 1056
rect 1069 944 1075 1016
rect 1101 984 1107 1336
rect 1149 1284 1155 1316
rect 1213 1284 1219 1476
rect 1229 1464 1235 1476
rect 1229 1324 1235 1336
rect 1373 1324 1379 1496
rect 1389 1404 1395 1496
rect 1533 1424 1539 1476
rect 1565 1464 1571 1616
rect 1565 1364 1571 1456
rect 1277 1304 1283 1316
rect 1117 1024 1123 1056
rect 1117 944 1123 1016
rect 1053 903 1059 916
rect 1044 897 1059 903
rect 989 704 995 856
rect 1021 717 1036 723
rect 1021 684 1027 717
rect 1069 704 1075 916
rect 1133 884 1139 1096
rect 1149 1084 1155 1276
rect 1165 1124 1171 1236
rect 1245 1164 1251 1296
rect 1229 1084 1235 1096
rect 1245 1084 1251 1156
rect 1101 704 1107 876
rect 1165 784 1171 916
rect 1181 784 1187 896
rect 1277 884 1283 1296
rect 1293 1144 1299 1236
rect 1309 1124 1315 1136
rect 1373 1084 1379 1156
rect 1421 1104 1427 1116
rect 1485 1104 1491 1336
rect 1549 1262 1555 1300
rect 1565 1244 1571 1356
rect 1581 1163 1587 1416
rect 1661 1384 1667 1737
rect 1693 1684 1699 1696
rect 1725 1544 1731 1876
rect 1757 1764 1763 1776
rect 1821 1744 1827 1796
rect 1837 1724 1843 1736
rect 1741 1524 1747 1716
rect 1853 1704 1859 1716
rect 1773 1564 1779 1636
rect 1805 1524 1811 1576
rect 1821 1524 1827 1556
rect 1837 1544 1843 1676
rect 1853 1664 1859 1676
rect 1741 1504 1747 1516
rect 1629 1304 1635 1316
rect 1597 1184 1603 1236
rect 1581 1157 1603 1163
rect 1389 1044 1395 1096
rect 1453 1084 1459 1096
rect 1405 1003 1411 1076
rect 1437 1024 1443 1076
rect 1485 1024 1491 1056
rect 1389 997 1411 1003
rect 1229 724 1235 736
rect 1037 684 1043 696
rect 1021 664 1027 676
rect 824 406 830 414
rect 838 406 844 414
rect 852 406 858 414
rect 866 406 872 414
rect 941 384 947 516
rect 653 324 659 376
rect 861 304 867 376
rect 1021 364 1027 556
rect 1053 544 1059 556
rect 461 144 467 276
rect 605 264 611 276
rect 541 184 547 236
rect 397 124 403 136
rect 493 124 499 156
rect 653 144 659 256
rect 781 244 787 256
rect 861 204 867 296
rect 877 244 883 356
rect 941 324 947 336
rect 1117 303 1123 696
rect 1133 657 1139 676
rect 1229 663 1235 696
rect 1245 663 1251 876
rect 1277 664 1283 716
rect 1325 704 1331 716
rect 1229 657 1251 663
rect 1229 564 1235 636
rect 1149 524 1155 536
rect 1149 444 1155 496
rect 1197 384 1203 516
rect 1245 464 1251 657
rect 1293 584 1299 676
rect 1325 664 1331 676
rect 1357 544 1363 956
rect 1389 944 1395 997
rect 1533 944 1539 1016
rect 1453 862 1459 900
rect 1405 657 1420 663
rect 1389 564 1395 656
rect 1405 584 1411 657
rect 1437 564 1443 716
rect 1533 704 1539 916
rect 1549 904 1555 916
rect 1581 904 1587 1036
rect 1597 984 1603 1157
rect 1629 1144 1635 1296
rect 1629 924 1635 956
rect 1693 924 1699 1216
rect 1725 1064 1731 1076
rect 1581 864 1587 896
rect 1597 884 1603 896
rect 1709 884 1715 896
rect 1741 884 1747 1456
rect 1757 1384 1763 1476
rect 1821 1324 1827 1436
rect 1773 1304 1779 1316
rect 1789 1264 1795 1316
rect 1837 1284 1843 1536
rect 1885 1504 1891 1836
rect 1901 1744 1907 1756
rect 1997 1744 2003 1856
rect 2072 1806 2078 1814
rect 2086 1806 2092 1814
rect 2100 1806 2106 1814
rect 2114 1806 2120 1814
rect 2173 1804 2179 1856
rect 2029 1784 2035 1796
rect 1949 1724 1955 1736
rect 1965 1704 1971 1716
rect 2029 1704 2035 1756
rect 1949 1543 1955 1676
rect 1940 1537 1955 1543
rect 1965 1524 1971 1696
rect 1917 1504 1923 1516
rect 1885 1464 1891 1496
rect 1853 1303 1859 1376
rect 1885 1344 1891 1456
rect 1901 1384 1907 1476
rect 1876 1317 1891 1323
rect 1853 1297 1868 1303
rect 1773 1257 1788 1263
rect 1773 1184 1779 1257
rect 1885 1224 1891 1317
rect 1917 1184 1923 1456
rect 1933 1324 1939 1496
rect 1949 1324 1955 1336
rect 1933 1124 1939 1316
rect 1965 1184 1971 1496
rect 2045 1384 2051 1456
rect 2072 1406 2078 1414
rect 2086 1406 2092 1414
rect 2100 1406 2106 1414
rect 2114 1406 2120 1414
rect 2077 1344 2083 1376
rect 1981 1184 1987 1216
rect 1757 924 1763 1076
rect 1773 884 1779 956
rect 1805 884 1811 956
rect 1885 944 1891 956
rect 1917 924 1923 956
rect 1869 904 1875 916
rect 1549 804 1555 836
rect 1613 664 1619 756
rect 1645 684 1651 796
rect 1709 720 1715 758
rect 1357 464 1363 516
rect 1245 384 1251 456
rect 1165 323 1171 336
rect 1165 317 1180 323
rect 1108 297 1123 303
rect 877 164 883 236
rect 957 124 963 196
rect 1053 183 1059 256
rect 1053 177 1068 183
rect 1069 164 1075 176
rect 1101 144 1107 296
rect 1133 264 1139 316
rect 1236 277 1251 283
rect 1149 124 1155 176
rect 1165 164 1171 276
rect 1245 184 1251 277
rect 1293 204 1299 276
rect 1165 144 1171 156
rect 1181 124 1187 136
rect 45 44 51 96
rect 781 44 787 100
rect 1229 103 1235 156
rect 1220 97 1235 103
rect 824 6 830 14
rect 838 6 844 14
rect 852 6 858 14
rect 866 6 872 14
rect 1117 -17 1123 36
rect 237 -23 243 -17
rect 1117 -23 1139 -17
rect 1261 -23 1267 196
rect 1389 164 1395 176
rect 1405 163 1411 436
rect 1421 384 1427 536
rect 1453 524 1459 636
rect 1613 564 1619 656
rect 1613 544 1619 556
rect 1645 544 1651 556
rect 1709 462 1715 500
rect 1725 484 1731 836
rect 1805 784 1811 856
rect 1901 784 1907 896
rect 1933 864 1939 1116
rect 1949 1104 1955 1176
rect 2013 1104 2019 1176
rect 2125 1124 2131 1336
rect 2141 1304 2147 1776
rect 2189 1704 2195 1716
rect 2253 1464 2259 1796
rect 2269 1784 2275 1876
rect 2269 1704 2275 1716
rect 2285 1504 2291 1896
rect 2557 1884 2563 1896
rect 2461 1864 2467 1876
rect 2573 1864 2579 1876
rect 2557 1857 2572 1863
rect 2397 1824 2403 1856
rect 2429 1763 2435 1836
rect 2493 1784 2499 1836
rect 2429 1757 2451 1763
rect 2445 1744 2451 1757
rect 2429 1584 2435 1696
rect 2445 1563 2451 1716
rect 2349 1520 2355 1558
rect 2429 1557 2451 1563
rect 2397 1484 2403 1496
rect 2189 1304 2195 1356
rect 2221 1324 2227 1356
rect 2285 1337 2300 1343
rect 2141 1144 2147 1296
rect 2173 1104 2179 1236
rect 2237 1104 2243 1136
rect 2180 1097 2188 1103
rect 2285 1084 2291 1337
rect 2333 1304 2339 1356
rect 2413 1344 2419 1356
rect 2429 1324 2435 1557
rect 2461 1524 2467 1716
rect 2477 1524 2483 1676
rect 2509 1564 2515 1636
rect 2461 1504 2467 1516
rect 2477 1364 2483 1516
rect 2349 1264 2355 1316
rect 2429 1124 2435 1316
rect 2461 1264 2467 1296
rect 2493 1283 2499 1316
rect 2509 1284 2515 1536
rect 2525 1523 2531 1836
rect 2557 1684 2563 1857
rect 2541 1544 2547 1676
rect 2573 1584 2579 1816
rect 2589 1784 2595 1896
rect 2749 1764 2755 1856
rect 2781 1844 2787 1876
rect 2525 1517 2547 1523
rect 2477 1277 2499 1283
rect 2461 1104 2467 1116
rect 2445 1084 2451 1096
rect 2045 984 2051 1036
rect 2072 1006 2078 1014
rect 2086 1006 2092 1014
rect 2100 1006 2106 1014
rect 2114 1006 2120 1014
rect 2157 984 2163 1056
rect 2173 1044 2179 1076
rect 1981 906 1987 956
rect 2029 944 2035 956
rect 2045 904 2051 956
rect 1981 744 1987 898
rect 2141 884 2147 956
rect 2173 924 2179 1036
rect 2189 944 2195 956
rect 2180 917 2188 923
rect 2157 884 2163 916
rect 2180 897 2195 903
rect 1741 524 1747 696
rect 1837 584 1843 676
rect 1885 664 1891 716
rect 1949 664 1955 736
rect 1981 704 1987 736
rect 1997 684 2003 696
rect 1517 320 1523 358
rect 1581 284 1587 416
rect 1773 384 1779 576
rect 1901 544 1907 636
rect 1789 524 1795 536
rect 1917 523 1923 576
rect 1997 564 2003 636
rect 2013 543 2019 716
rect 2093 704 2099 876
rect 2189 844 2195 897
rect 2189 744 2195 836
rect 2205 744 2211 1036
rect 2285 904 2291 936
rect 2317 904 2323 956
rect 2333 924 2339 1016
rect 2413 964 2419 1036
rect 2429 924 2435 1036
rect 2461 964 2467 1096
rect 2477 1044 2483 1277
rect 2509 1144 2515 1276
rect 2525 1144 2531 1436
rect 2541 1344 2547 1517
rect 2557 1324 2563 1556
rect 2573 1124 2579 1436
rect 2589 1404 2595 1636
rect 2605 1383 2611 1736
rect 2749 1643 2755 1756
rect 2861 1724 2867 1896
rect 2845 1662 2851 1700
rect 2733 1637 2755 1643
rect 2653 1484 2659 1496
rect 2596 1377 2611 1383
rect 2653 1324 2659 1476
rect 2733 1464 2739 1637
rect 2829 1520 2835 1558
rect 2861 1504 2867 1716
rect 2733 1404 2739 1456
rect 2781 1364 2787 1396
rect 2589 1304 2595 1316
rect 2877 1244 2883 1300
rect 2509 1104 2515 1116
rect 2525 1044 2531 1096
rect 2532 1037 2547 1043
rect 2509 944 2515 956
rect 2541 924 2547 1037
rect 2093 684 2099 696
rect 2141 684 2147 696
rect 2072 606 2078 614
rect 2086 606 2092 614
rect 2100 606 2106 614
rect 2114 606 2120 614
rect 2141 544 2147 636
rect 2157 544 2163 716
rect 2189 544 2195 556
rect 2013 537 2035 543
rect 1901 517 1923 523
rect 1837 464 1843 516
rect 1837 324 1843 376
rect 1853 304 1859 516
rect 1885 504 1891 516
rect 1901 504 1907 517
rect 1917 464 1923 496
rect 1933 424 1939 516
rect 1949 444 1955 516
rect 1965 464 1971 536
rect 2013 497 2019 516
rect 2029 504 2035 537
rect 2221 543 2227 856
rect 2269 704 2275 896
rect 2461 864 2467 896
rect 2317 704 2323 736
rect 2301 683 2307 696
rect 2301 677 2316 683
rect 2237 584 2243 656
rect 2365 624 2371 656
rect 2301 564 2307 576
rect 2221 537 2236 543
rect 2157 504 2163 536
rect 2189 524 2195 536
rect 1613 204 1619 256
rect 1565 164 1571 196
rect 1396 157 1411 163
rect 1277 144 1283 156
rect 1293 124 1299 136
rect 1693 124 1699 296
rect 1933 284 1939 396
rect 2077 384 2083 496
rect 2125 404 2131 436
rect 2157 324 2163 496
rect 2157 284 2163 316
rect 1853 184 1859 256
rect 2045 164 2051 256
rect 2072 206 2078 214
rect 2086 206 2092 214
rect 2100 206 2106 214
rect 2114 206 2120 214
rect 2205 184 2211 256
rect 2221 184 2227 537
rect 2237 324 2243 376
rect 2253 344 2259 556
rect 2381 544 2387 676
rect 2397 524 2403 696
rect 2413 544 2419 556
rect 2445 524 2451 676
rect 2461 544 2467 696
rect 2301 324 2307 356
rect 2365 304 2371 336
rect 2381 324 2387 416
rect 2253 284 2259 296
rect 2285 144 2291 276
rect 2301 184 2307 276
rect 2381 264 2387 316
rect 2397 304 2403 496
rect 2477 484 2483 876
rect 2525 844 2531 896
rect 2541 723 2547 836
rect 2621 784 2627 836
rect 2541 717 2556 723
rect 2573 563 2579 636
rect 2637 603 2643 1136
rect 2845 1120 2851 1158
rect 2669 1064 2675 1096
rect 2749 1023 2755 1056
rect 2749 1017 2771 1023
rect 2765 964 2771 1017
rect 2765 843 2771 956
rect 2877 924 2883 1096
rect 2861 862 2867 900
rect 2765 837 2787 843
rect 2781 764 2787 837
rect 2781 664 2787 756
rect 2877 704 2883 916
rect 2909 724 2915 776
rect 2621 597 2643 603
rect 2564 557 2579 563
rect 2557 544 2563 556
rect 2589 524 2595 576
rect 2477 444 2483 476
rect 2573 464 2579 496
rect 2605 484 2611 516
rect 2413 344 2419 436
rect 2477 324 2483 396
rect 2493 344 2499 436
rect 2509 384 2515 436
rect 2493 324 2499 336
rect 2541 324 2547 376
rect 2573 323 2579 456
rect 2589 404 2595 436
rect 2573 317 2595 323
rect 2445 284 2451 316
rect 2557 304 2563 316
rect 2493 284 2499 296
rect 2589 284 2595 317
rect 2589 264 2595 276
rect 2461 164 2467 256
rect 2541 204 2547 236
rect 2493 144 2499 196
rect 1277 104 1283 116
rect 1661 62 1667 100
rect 1741 -23 1747 136
rect 2589 124 2595 196
rect 2621 124 2627 597
rect 2829 584 2835 616
rect 2877 584 2883 696
rect 2637 504 2643 576
rect 2653 524 2659 536
rect 2749 524 2755 536
rect 2669 484 2675 516
rect 2701 424 2707 516
rect 2717 464 2723 516
rect 2765 504 2771 516
rect 2781 504 2787 516
rect 2829 504 2835 536
rect 2781 384 2787 436
rect 2637 324 2643 376
rect 2637 204 2643 296
rect 2653 184 2659 356
rect 2845 304 2851 576
rect 2877 544 2883 556
rect 2861 324 2867 516
rect 2685 184 2691 216
rect 2861 184 2867 276
rect 2717 124 2723 176
rect 2740 137 2755 143
rect 2685 104 2691 116
rect 2749 104 2755 137
rect 2765 124 2771 156
rect 2813 144 2819 176
rect 2877 104 2883 536
rect 2893 124 2899 496
rect 1917 44 1923 96
rect 2557 44 2563 100
rect 2781 84 2787 96
rect 2765 64 2771 76
rect 2893 64 2899 96
rect 2909 84 2915 476
rect 2925 384 2931 556
rect 2941 124 2947 436
<< m3contact >>
rect 12 1936 20 1944
rect 28 1936 36 1944
rect 284 1936 292 1944
rect 300 1936 308 1944
rect 332 1936 340 1944
rect 92 1916 100 1924
rect 204 1916 212 1924
rect 60 1896 68 1904
rect 140 1896 148 1904
rect 60 1876 68 1884
rect 140 1876 148 1884
rect 12 1856 20 1864
rect 108 1856 116 1864
rect 44 1776 52 1784
rect 44 1756 52 1764
rect 92 1756 100 1764
rect 60 1736 68 1744
rect 92 1736 100 1744
rect 12 1696 20 1704
rect 28 1696 36 1704
rect 220 1876 228 1884
rect 316 1916 324 1924
rect 380 1916 388 1924
rect 460 1916 468 1924
rect 364 1896 372 1904
rect 188 1856 196 1864
rect 252 1856 260 1864
rect 268 1856 276 1864
rect 348 1856 356 1864
rect 204 1796 212 1804
rect 316 1796 324 1804
rect 188 1756 196 1764
rect 300 1756 308 1764
rect 172 1736 180 1744
rect 156 1716 164 1724
rect 76 1676 84 1684
rect 108 1556 116 1564
rect 44 1516 52 1524
rect 92 1516 100 1524
rect 236 1716 244 1724
rect 252 1716 260 1724
rect 140 1696 148 1704
rect 204 1696 212 1704
rect 252 1696 260 1704
rect 332 1756 340 1764
rect 348 1716 356 1724
rect 364 1716 372 1724
rect 444 1896 452 1904
rect 588 1916 596 1924
rect 556 1896 564 1904
rect 428 1856 436 1864
rect 476 1796 484 1804
rect 476 1756 484 1764
rect 508 1756 516 1764
rect 396 1736 404 1744
rect 268 1656 276 1664
rect 204 1516 212 1524
rect 332 1576 340 1584
rect 316 1536 324 1544
rect 140 1496 148 1504
rect 172 1496 180 1504
rect 204 1496 212 1504
rect 236 1496 244 1504
rect 284 1496 292 1504
rect 348 1496 356 1504
rect 12 1456 20 1464
rect 252 1476 260 1484
rect 284 1476 292 1484
rect 412 1716 420 1724
rect 428 1696 436 1704
rect 830 2006 838 2014
rect 844 2006 852 2014
rect 858 2006 866 2014
rect 684 1916 692 1924
rect 636 1896 644 1904
rect 716 1896 724 1904
rect 908 1816 916 1824
rect 764 1796 772 1804
rect 748 1776 756 1784
rect 572 1756 580 1764
rect 748 1736 756 1744
rect 972 1736 980 1744
rect 604 1716 612 1724
rect 860 1716 868 1724
rect 1036 1716 1044 1724
rect 460 1676 468 1684
rect 412 1576 420 1584
rect 428 1536 436 1544
rect 588 1676 596 1684
rect 524 1536 532 1544
rect 652 1696 660 1704
rect 908 1696 916 1704
rect 956 1696 964 1704
rect 620 1656 628 1664
rect 604 1556 612 1564
rect 444 1516 452 1524
rect 540 1516 548 1524
rect 76 1456 84 1464
rect 316 1456 324 1464
rect 460 1456 468 1464
rect 204 1436 212 1444
rect 316 1396 324 1404
rect 300 1376 308 1384
rect 172 1356 180 1364
rect 268 1356 276 1364
rect 44 1316 52 1324
rect 108 1316 114 1324
rect 114 1316 116 1324
rect 12 1296 20 1304
rect 140 1196 148 1204
rect 364 1356 372 1364
rect 380 1336 388 1344
rect 332 1176 340 1184
rect 252 1096 260 1104
rect 380 1096 388 1104
rect 140 936 148 944
rect 140 676 148 684
rect 364 956 372 964
rect 348 936 356 944
rect 444 1396 452 1404
rect 476 1376 484 1384
rect 604 1456 612 1464
rect 556 1396 564 1404
rect 556 1356 564 1364
rect 572 1356 580 1364
rect 460 1336 468 1344
rect 492 1336 500 1344
rect 636 1456 644 1464
rect 830 1606 838 1614
rect 844 1606 852 1614
rect 858 1606 866 1614
rect 732 1536 740 1544
rect 876 1536 884 1544
rect 780 1516 788 1524
rect 924 1516 932 1524
rect 764 1496 772 1504
rect 956 1496 964 1504
rect 748 1476 756 1484
rect 924 1476 932 1484
rect 812 1456 820 1464
rect 1004 1456 1012 1464
rect 700 1436 708 1444
rect 892 1436 900 1444
rect 652 1396 660 1404
rect 716 1356 724 1364
rect 748 1356 756 1364
rect 508 1316 516 1324
rect 620 1316 628 1324
rect 828 1316 836 1324
rect 716 1276 724 1284
rect 830 1206 838 1214
rect 844 1206 852 1214
rect 858 1206 866 1214
rect 556 1196 564 1204
rect 908 1136 916 1144
rect 684 1116 692 1124
rect 764 1116 772 1124
rect 812 1116 820 1124
rect 492 1076 500 1084
rect 524 1036 532 1044
rect 492 1016 500 1024
rect 556 996 564 1004
rect 556 956 564 964
rect 444 916 452 924
rect 428 876 436 884
rect 332 856 340 864
rect 412 856 420 864
rect 332 716 340 724
rect 412 716 420 724
rect 476 876 484 884
rect 524 876 532 884
rect 588 776 596 784
rect 348 676 356 684
rect 172 656 180 664
rect 140 536 148 544
rect 140 276 148 284
rect 348 536 356 544
rect 460 676 468 684
rect 508 676 516 684
rect 572 676 580 684
rect 508 656 516 664
rect 492 576 500 584
rect 444 516 452 524
rect 364 496 372 504
rect 332 456 340 464
rect 332 316 340 324
rect 252 296 260 304
rect 172 236 180 244
rect 140 136 148 144
rect 348 276 356 284
rect 396 456 404 464
rect 428 476 436 484
rect 412 316 420 324
rect 476 476 484 484
rect 796 1096 804 1104
rect 700 1076 708 1084
rect 764 1036 772 1044
rect 716 996 724 1004
rect 956 1116 964 1124
rect 1228 1996 1236 2004
rect 1276 1996 1284 2004
rect 1100 1916 1108 1924
rect 2348 1916 2356 1924
rect 2412 1916 2420 1924
rect 1180 1896 1188 1904
rect 1260 1896 1266 1904
rect 1266 1896 1268 1904
rect 1836 1896 1844 1904
rect 2092 1896 2100 1904
rect 2556 1896 2564 1904
rect 2588 1896 2596 1904
rect 1132 1876 1140 1884
rect 1132 1856 1140 1864
rect 1164 1816 1172 1824
rect 1084 1696 1092 1704
rect 1148 1636 1156 1644
rect 1452 1856 1460 1864
rect 1420 1816 1428 1824
rect 1500 1816 1508 1824
rect 1468 1736 1476 1744
rect 1292 1716 1300 1724
rect 1340 1716 1348 1724
rect 1372 1716 1380 1724
rect 1196 1616 1204 1624
rect 1244 1616 1252 1624
rect 1100 1536 1108 1544
rect 1164 1536 1172 1544
rect 1196 1536 1204 1544
rect 1068 1516 1076 1524
rect 1132 1516 1140 1524
rect 1244 1516 1252 1524
rect 1084 1476 1092 1484
rect 1084 1456 1092 1464
rect 1116 1456 1124 1464
rect 1068 1436 1076 1444
rect 1020 1336 1028 1344
rect 1068 1336 1076 1344
rect 1116 1336 1124 1344
rect 1148 1496 1156 1504
rect 2204 1876 2212 1884
rect 2268 1876 2276 1884
rect 1500 1616 1508 1624
rect 1564 1616 1572 1624
rect 1324 1496 1332 1504
rect 1372 1496 1380 1504
rect 1436 1496 1444 1504
rect 1292 1476 1300 1484
rect 1052 1296 1060 1304
rect 1084 1276 1092 1284
rect 1020 1116 1028 1124
rect 988 1096 996 1104
rect 1036 1096 1044 1104
rect 1052 1096 1060 1104
rect 812 1016 820 1024
rect 732 936 740 944
rect 844 896 852 904
rect 700 816 708 824
rect 764 816 772 824
rect 668 696 676 704
rect 830 806 838 814
rect 844 806 852 814
rect 858 806 866 814
rect 876 696 884 704
rect 860 676 862 684
rect 862 676 868 684
rect 700 656 708 664
rect 748 576 756 584
rect 780 576 788 584
rect 588 556 596 564
rect 684 556 692 564
rect 716 556 724 564
rect 556 536 564 544
rect 620 536 628 544
rect 588 516 596 524
rect 636 516 644 524
rect 700 516 708 524
rect 828 536 836 544
rect 764 516 772 524
rect 1068 1056 1076 1064
rect 1068 1016 1076 1024
rect 1132 1296 1140 1304
rect 1196 1296 1204 1304
rect 1228 1456 1236 1464
rect 1532 1416 1540 1424
rect 1388 1396 1396 1404
rect 1580 1416 1588 1424
rect 1452 1356 1460 1364
rect 1564 1356 1572 1364
rect 1228 1316 1236 1324
rect 1372 1316 1380 1324
rect 1244 1296 1252 1304
rect 1276 1296 1284 1304
rect 1148 1276 1156 1284
rect 1212 1276 1220 1284
rect 1116 1016 1124 1024
rect 1100 976 1108 984
rect 1084 936 1092 944
rect 1036 916 1044 924
rect 1068 916 1076 924
rect 988 856 996 864
rect 1004 736 1012 744
rect 972 696 980 704
rect 1244 1156 1252 1164
rect 1164 1116 1172 1124
rect 1196 1116 1204 1124
rect 1228 1116 1236 1124
rect 1260 1096 1268 1104
rect 1148 1076 1156 1084
rect 1180 1076 1188 1084
rect 1228 1076 1236 1084
rect 1260 1076 1268 1084
rect 1196 976 1204 984
rect 1100 876 1108 884
rect 1132 876 1140 884
rect 1180 896 1188 904
rect 1372 1156 1380 1164
rect 1292 1136 1300 1144
rect 1308 1136 1316 1144
rect 1356 1096 1364 1104
rect 1420 1116 1428 1124
rect 1564 1236 1572 1244
rect 1516 1176 1524 1184
rect 1676 1736 1684 1744
rect 1676 1716 1684 1724
rect 1692 1676 1700 1684
rect 1756 1856 1764 1864
rect 2172 1856 2180 1864
rect 1884 1836 1892 1844
rect 1916 1836 1924 1844
rect 1820 1796 1828 1804
rect 1756 1776 1764 1784
rect 1740 1736 1748 1744
rect 1788 1736 1796 1744
rect 1836 1736 1844 1744
rect 1836 1716 1844 1724
rect 1724 1536 1732 1544
rect 1852 1696 1860 1704
rect 1852 1676 1860 1684
rect 1804 1576 1812 1584
rect 1772 1556 1780 1564
rect 1772 1536 1780 1544
rect 1820 1556 1828 1564
rect 1836 1536 1844 1544
rect 1740 1516 1748 1524
rect 1772 1496 1780 1504
rect 1724 1356 1732 1364
rect 1692 1336 1700 1344
rect 1628 1296 1636 1304
rect 1724 1296 1732 1304
rect 1596 1236 1604 1244
rect 1324 1076 1332 1084
rect 1324 1056 1332 1064
rect 1356 1056 1364 1064
rect 1452 1076 1460 1084
rect 1388 1036 1396 1044
rect 1580 1036 1588 1044
rect 1436 1016 1444 1024
rect 1484 1016 1492 1024
rect 1532 1016 1540 1024
rect 1244 876 1252 884
rect 1276 876 1284 884
rect 1164 776 1172 784
rect 1228 736 1236 744
rect 1036 696 1044 704
rect 1068 696 1076 704
rect 1116 696 1124 704
rect 1020 676 1028 684
rect 1084 676 1092 684
rect 924 576 932 584
rect 1052 556 1060 564
rect 652 496 660 504
rect 732 496 740 504
rect 908 496 916 504
rect 830 406 838 414
rect 844 406 852 414
rect 858 406 866 414
rect 860 376 868 384
rect 940 376 948 384
rect 508 316 516 324
rect 876 356 884 364
rect 1020 356 1028 364
rect 636 296 644 304
rect 748 276 756 284
rect 444 156 452 164
rect 604 256 612 264
rect 652 256 660 264
rect 540 236 548 244
rect 492 156 500 164
rect 348 136 356 144
rect 396 136 404 144
rect 444 136 452 144
rect 460 136 468 144
rect 780 236 788 244
rect 940 316 948 324
rect 1068 316 1076 324
rect 1020 296 1028 304
rect 1052 296 1060 304
rect 1132 676 1140 684
rect 1276 716 1284 724
rect 1324 716 1332 724
rect 1340 696 1348 704
rect 1292 676 1300 684
rect 1148 536 1156 544
rect 1324 656 1332 664
rect 1484 916 1492 924
rect 1532 916 1540 924
rect 1452 776 1460 784
rect 1372 716 1380 724
rect 1436 716 1444 724
rect 1692 1216 1700 1224
rect 1628 1136 1636 1144
rect 1628 956 1636 964
rect 1644 936 1652 944
rect 1708 1076 1716 1084
rect 1724 1056 1732 1064
rect 1548 896 1556 904
rect 1676 896 1684 904
rect 1772 1316 1780 1324
rect 1820 1316 1828 1324
rect 1916 1756 1924 1764
rect 2078 1806 2086 1814
rect 2092 1806 2100 1814
rect 2106 1806 2114 1814
rect 2028 1796 2036 1804
rect 2172 1796 2180 1804
rect 2252 1796 2260 1804
rect 2140 1776 2148 1784
rect 2172 1776 2180 1784
rect 2028 1756 2036 1764
rect 1900 1736 1908 1744
rect 2012 1736 2020 1744
rect 1948 1716 1956 1724
rect 2076 1736 2084 1744
rect 1964 1696 1972 1704
rect 1916 1576 1924 1584
rect 1932 1536 1940 1544
rect 1916 1516 1924 1524
rect 1964 1516 1972 1524
rect 1996 1516 2004 1524
rect 1932 1496 1940 1504
rect 1900 1476 1908 1484
rect 1852 1376 1860 1384
rect 1916 1456 1924 1464
rect 1884 1336 1892 1344
rect 1820 1276 1828 1284
rect 1836 1276 1844 1284
rect 1852 1276 1860 1284
rect 1788 1256 1796 1264
rect 1884 1216 1892 1224
rect 1948 1316 1956 1324
rect 2078 1406 2086 1414
rect 2092 1406 2100 1414
rect 2106 1406 2114 1414
rect 2044 1376 2052 1384
rect 2076 1376 2084 1384
rect 1996 1356 2004 1364
rect 2124 1336 2132 1344
rect 2028 1316 2036 1324
rect 1980 1216 1988 1224
rect 1948 1176 1956 1184
rect 1964 1176 1972 1184
rect 2012 1176 2020 1184
rect 1932 1116 1940 1124
rect 1804 1076 1812 1084
rect 1884 956 1892 964
rect 1916 956 1924 964
rect 1788 936 1796 944
rect 1820 916 1828 924
rect 1916 916 1924 924
rect 1868 896 1876 904
rect 1916 896 1924 904
rect 1596 876 1604 884
rect 1660 876 1668 884
rect 1708 876 1716 884
rect 1740 876 1748 884
rect 1772 876 1780 884
rect 1804 876 1812 884
rect 1580 856 1588 864
rect 1804 856 1812 864
rect 1548 796 1556 804
rect 1644 796 1652 804
rect 1612 756 1620 764
rect 1388 556 1396 564
rect 1308 536 1316 544
rect 1356 536 1364 544
rect 1420 536 1428 544
rect 1260 516 1268 524
rect 1372 516 1380 524
rect 1244 456 1252 464
rect 1356 456 1364 464
rect 1132 316 1140 324
rect 956 276 964 284
rect 876 236 884 244
rect 860 196 868 204
rect 956 196 964 204
rect 508 136 516 144
rect 844 136 852 144
rect 1068 176 1076 184
rect 1116 276 1124 284
rect 1164 296 1172 304
rect 1164 276 1172 284
rect 1148 176 1156 184
rect 1052 136 1060 144
rect 1100 136 1108 144
rect 1308 276 1316 284
rect 1260 196 1268 204
rect 1292 196 1300 204
rect 1164 156 1172 164
rect 1180 136 1188 144
rect 332 116 334 124
rect 334 116 340 124
rect 444 116 452 124
rect 1100 116 1108 124
rect 1196 116 1204 124
rect 1036 96 1044 104
rect 1212 96 1220 104
rect 830 6 838 14
rect 844 6 852 14
rect 858 6 866 14
rect 1388 176 1396 184
rect 1276 156 1284 164
rect 1644 556 1652 564
rect 1612 536 1620 544
rect 1452 516 1460 524
rect 2156 1756 2164 1764
rect 2188 1696 2196 1704
rect 2268 1716 2276 1724
rect 2380 1876 2388 1884
rect 2572 1876 2580 1884
rect 2460 1856 2468 1864
rect 2492 1836 2500 1844
rect 2396 1816 2404 1824
rect 2332 1736 2340 1744
rect 2428 1736 2436 1744
rect 2300 1716 2308 1724
rect 2444 1716 2452 1724
rect 2460 1716 2468 1724
rect 2428 1696 2436 1704
rect 2284 1476 2292 1484
rect 2396 1476 2404 1484
rect 2252 1456 2260 1464
rect 2220 1356 2228 1364
rect 2284 1356 2292 1364
rect 2412 1356 2420 1364
rect 2156 1336 2164 1344
rect 2204 1336 2212 1344
rect 2140 1296 2148 1304
rect 2188 1296 2196 1304
rect 2252 1296 2260 1304
rect 2236 1136 2244 1144
rect 2140 1096 2148 1104
rect 2172 1096 2180 1104
rect 2444 1536 2452 1544
rect 2492 1696 2500 1704
rect 2476 1676 2484 1684
rect 2508 1556 2516 1564
rect 2508 1536 2516 1544
rect 2460 1516 2468 1524
rect 2460 1496 2468 1504
rect 2476 1356 2484 1364
rect 2460 1336 2468 1344
rect 2428 1316 2436 1324
rect 2300 1296 2308 1304
rect 2332 1296 2340 1304
rect 2380 1276 2388 1284
rect 2348 1256 2356 1264
rect 2476 1296 2484 1304
rect 2540 1716 2548 1724
rect 2572 1816 2580 1824
rect 2556 1676 2564 1684
rect 2780 1836 2788 1844
rect 2604 1736 2612 1744
rect 2556 1556 2564 1564
rect 2524 1496 2532 1504
rect 2460 1256 2468 1264
rect 2428 1116 2436 1124
rect 2460 1116 2468 1124
rect 2396 1096 2404 1104
rect 2444 1096 2452 1104
rect 2172 1076 2180 1084
rect 2284 1076 2292 1084
rect 2300 1076 2308 1084
rect 2428 1076 2436 1084
rect 2156 1056 2164 1064
rect 1980 1036 1988 1044
rect 2078 1006 2086 1014
rect 2092 1006 2100 1014
rect 2106 1006 2114 1014
rect 2220 1056 2228 1064
rect 2268 1056 2276 1064
rect 2428 1036 2436 1044
rect 2044 976 2052 984
rect 1980 956 1988 964
rect 2028 956 2036 964
rect 2140 956 2148 964
rect 1964 936 1972 944
rect 2028 916 2036 924
rect 1932 856 1940 864
rect 2044 896 2052 904
rect 2188 956 2196 964
rect 2172 916 2180 924
rect 2092 876 2100 884
rect 2156 876 2164 884
rect 1948 736 1956 744
rect 1820 716 1828 724
rect 1852 716 1860 724
rect 1852 696 1860 704
rect 1788 676 1796 684
rect 1820 676 1828 684
rect 1916 696 1924 704
rect 1916 676 1924 684
rect 2012 716 2020 724
rect 1980 696 1988 704
rect 1996 676 2004 684
rect 1884 656 1892 664
rect 1772 576 1780 584
rect 1836 576 1844 584
rect 1740 516 1748 524
rect 1724 476 1732 484
rect 1580 416 1588 424
rect 1916 576 1924 584
rect 1900 536 1908 544
rect 1788 516 1796 524
rect 1852 516 1860 524
rect 1996 556 2004 564
rect 2188 836 2196 844
rect 2332 1016 2340 1024
rect 2284 936 2292 944
rect 2268 916 2276 924
rect 2412 956 2420 964
rect 2508 1276 2516 1284
rect 2492 1256 2500 1264
rect 2540 1316 2548 1324
rect 2556 1316 2564 1324
rect 2524 1136 2532 1144
rect 2588 1396 2596 1404
rect 2780 1736 2788 1744
rect 2652 1476 2660 1484
rect 2764 1476 2772 1484
rect 2732 1456 2740 1464
rect 2732 1396 2740 1404
rect 2780 1396 2788 1404
rect 2812 1336 2820 1344
rect 2588 1316 2596 1324
rect 2652 1316 2660 1324
rect 2700 1316 2708 1324
rect 2620 1296 2628 1304
rect 2636 1136 2644 1144
rect 2492 1116 2500 1124
rect 2556 1116 2564 1124
rect 2572 1116 2580 1124
rect 2508 1096 2516 1104
rect 2588 1096 2594 1104
rect 2594 1096 2596 1104
rect 2492 1076 2500 1084
rect 2476 1036 2484 1044
rect 2524 1036 2532 1044
rect 2460 956 2468 964
rect 2508 956 2516 964
rect 2476 936 2484 944
rect 2492 916 2500 924
rect 2236 896 2244 904
rect 2268 896 2276 904
rect 2300 896 2308 904
rect 2316 896 2324 904
rect 2444 896 2452 904
rect 2604 896 2612 904
rect 2220 856 2228 864
rect 2156 736 2164 744
rect 2204 736 2212 744
rect 2156 716 2164 724
rect 2028 696 2036 704
rect 2140 696 2148 704
rect 2044 676 2052 684
rect 2092 676 2100 684
rect 2060 636 2068 644
rect 2140 636 2148 644
rect 2078 606 2086 614
rect 2092 606 2100 614
rect 2106 606 2114 614
rect 2204 696 2212 704
rect 2188 556 2196 564
rect 1836 456 1844 464
rect 1884 496 1892 504
rect 1868 476 1876 484
rect 1884 456 1892 464
rect 1916 456 1924 464
rect 2012 516 2020 524
rect 2156 536 2164 544
rect 2364 876 2372 884
rect 2412 876 2420 884
rect 2476 876 2484 884
rect 2428 856 2436 864
rect 2460 856 2468 864
rect 2316 736 2324 744
rect 2428 716 2436 724
rect 2428 696 2436 704
rect 2348 656 2356 664
rect 2364 616 2372 624
rect 2236 576 2244 584
rect 2300 576 2308 584
rect 2284 556 2292 564
rect 2332 556 2340 564
rect 2188 516 2196 524
rect 1996 476 2004 484
rect 1964 456 1972 464
rect 1948 436 1956 444
rect 1932 416 1940 424
rect 1932 396 1940 404
rect 1692 296 1700 304
rect 1852 296 1860 304
rect 1612 256 1620 264
rect 1564 196 1572 204
rect 1612 196 1620 204
rect 1292 136 1300 144
rect 1388 136 1396 144
rect 1596 136 1604 144
rect 2124 396 2132 404
rect 2076 376 2084 384
rect 2124 376 2132 384
rect 2204 436 2212 444
rect 2156 316 2164 324
rect 1852 256 1860 264
rect 1964 256 1972 264
rect 2044 256 2052 264
rect 2204 256 2212 264
rect 2078 206 2086 214
rect 2092 206 2100 214
rect 2106 206 2114 214
rect 2236 376 2244 384
rect 2316 536 2324 544
rect 2412 536 2420 544
rect 2428 536 2436 544
rect 2460 536 2468 544
rect 2364 516 2372 524
rect 2396 496 2404 504
rect 2268 456 2276 464
rect 2380 416 2388 424
rect 2300 356 2308 364
rect 2252 336 2260 344
rect 2364 336 2372 344
rect 2252 296 2260 304
rect 2300 296 2308 304
rect 2300 276 2308 284
rect 2364 276 2372 284
rect 2220 176 2228 184
rect 2044 156 2052 164
rect 2556 876 2564 884
rect 2524 836 2532 844
rect 2620 836 2628 844
rect 2524 696 2532 704
rect 2556 676 2564 684
rect 2780 1076 2788 1084
rect 2668 1056 2676 1064
rect 2796 936 2804 944
rect 2780 756 2788 764
rect 2812 676 2820 684
rect 2828 616 2836 624
rect 2588 576 2596 584
rect 2556 536 2564 544
rect 2524 516 2532 524
rect 2556 516 2564 524
rect 2604 516 2612 524
rect 2476 476 2484 484
rect 2572 456 2580 464
rect 2412 436 2420 444
rect 2476 436 2484 444
rect 2508 436 2516 444
rect 2476 396 2484 404
rect 2428 356 2436 364
rect 2508 376 2516 384
rect 2540 376 2548 384
rect 2492 336 2500 344
rect 2444 316 2452 324
rect 2492 316 2500 324
rect 2556 316 2564 324
rect 2588 396 2596 404
rect 2492 296 2500 304
rect 2572 296 2580 304
rect 2588 276 2596 284
rect 2316 256 2324 264
rect 2380 256 2388 264
rect 2460 256 2468 264
rect 2492 196 2500 204
rect 2540 196 2548 204
rect 2588 196 2596 204
rect 2460 156 2468 164
rect 1740 136 1748 144
rect 2012 136 2020 144
rect 2284 136 2292 144
rect 1276 96 1284 104
rect 1324 96 1332 104
rect 1404 96 1412 104
rect 2636 576 2644 584
rect 2844 576 2852 584
rect 2876 576 2884 584
rect 2652 536 2660 544
rect 2748 536 2756 544
rect 2828 536 2836 544
rect 2668 516 2676 524
rect 2716 516 2724 524
rect 2764 516 2772 524
rect 2652 436 2660 444
rect 2780 496 2788 504
rect 2796 476 2804 484
rect 2716 456 2724 464
rect 2700 416 2708 424
rect 2780 376 2788 384
rect 2652 356 2660 364
rect 2636 196 2644 204
rect 2876 556 2884 564
rect 2924 556 2932 564
rect 2892 536 2900 544
rect 2860 316 2868 324
rect 2732 276 2740 284
rect 2860 276 2868 284
rect 2764 256 2772 264
rect 2684 216 2692 224
rect 2716 176 2724 184
rect 2812 176 2820 184
rect 2636 136 2644 144
rect 2764 156 2772 164
rect 2732 136 2740 144
rect 2124 116 2132 124
rect 2380 116 2388 124
rect 2620 116 2628 124
rect 2684 116 2692 124
rect 2828 116 2836 124
rect 2892 496 2900 504
rect 2908 476 2916 484
rect 2668 96 2676 104
rect 2780 96 2788 104
rect 2860 96 2868 104
rect 2892 96 2900 104
rect 2764 76 2772 84
rect 2940 116 2948 124
<< metal3 >>
rect 824 2014 872 2016
rect 824 2006 828 2014
rect 838 2006 844 2014
rect 852 2006 858 2014
rect 868 2006 872 2014
rect 824 2004 872 2006
rect 1236 1997 1276 2003
rect -19 1937 12 1943
rect 36 1937 284 1943
rect 308 1937 332 1943
rect 100 1917 204 1923
rect 324 1917 380 1923
rect 388 1917 460 1923
rect 596 1917 684 1923
rect 692 1917 1100 1923
rect 2356 1917 2412 1923
rect -19 1897 60 1903
rect 116 1897 140 1903
rect 308 1897 364 1903
rect 452 1897 556 1903
rect 564 1897 636 1903
rect 644 1897 716 1903
rect 1188 1897 1260 1903
rect 1844 1897 2092 1903
rect 2564 1897 2588 1903
rect 68 1877 140 1883
rect 228 1877 355 1883
rect 349 1864 355 1877
rect 2212 1877 2268 1883
rect 2388 1877 2572 1883
rect 20 1857 108 1863
rect 116 1857 188 1863
rect 260 1857 268 1863
rect 276 1857 300 1863
rect 356 1857 428 1863
rect 1140 1857 1452 1863
rect 1764 1857 2172 1863
rect 2468 1857 2508 1863
rect 1892 1837 1916 1843
rect 2500 1837 2780 1843
rect 788 1817 908 1823
rect 916 1817 1164 1823
rect 1172 1817 1420 1823
rect 1428 1817 1500 1823
rect 2404 1817 2572 1823
rect 2072 1814 2120 1816
rect 2072 1806 2076 1814
rect 2086 1806 2092 1814
rect 2100 1806 2106 1814
rect 2116 1806 2120 1814
rect 2072 1804 2120 1806
rect 212 1797 316 1803
rect 484 1797 764 1803
rect 1828 1797 2028 1803
rect 2180 1797 2252 1803
rect 52 1777 748 1783
rect 1764 1777 2140 1783
rect 2148 1777 2172 1783
rect 52 1757 92 1763
rect 196 1757 300 1763
rect 340 1757 476 1763
rect 516 1757 572 1763
rect 1924 1757 2028 1763
rect 2036 1757 2156 1763
rect 68 1737 92 1743
rect 180 1737 396 1743
rect 404 1737 748 1743
rect 756 1737 972 1743
rect 1476 1737 1676 1743
rect 1748 1737 1788 1743
rect 1844 1737 1900 1743
rect 2020 1737 2076 1743
rect 2084 1737 2332 1743
rect 2388 1737 2428 1743
rect 2612 1737 2780 1743
rect 164 1717 236 1723
rect 260 1717 348 1723
rect 372 1717 412 1723
rect 612 1717 860 1723
rect 1044 1717 1292 1723
rect 1300 1717 1340 1723
rect 1348 1717 1372 1723
rect 1684 1717 1836 1723
rect 1956 1717 2268 1723
rect 2308 1717 2444 1723
rect 2468 1717 2540 1723
rect -19 1697 12 1703
rect 36 1697 140 1703
rect 148 1697 204 1703
rect 212 1697 252 1703
rect 436 1697 652 1703
rect 916 1697 956 1703
rect 964 1697 1084 1703
rect 1860 1697 1964 1703
rect 2196 1697 2380 1703
rect 2436 1697 2492 1703
rect 84 1677 460 1683
rect 468 1677 588 1683
rect 1700 1677 1852 1683
rect 2484 1677 2556 1683
rect 276 1657 620 1663
rect 1140 1637 1148 1643
rect 1204 1617 1244 1623
rect 1508 1617 1564 1623
rect 824 1614 872 1616
rect 824 1606 828 1614
rect 838 1606 844 1614
rect 852 1606 858 1614
rect 868 1606 872 1614
rect 824 1604 872 1606
rect 340 1577 412 1583
rect 1812 1577 1916 1583
rect 116 1557 604 1563
rect 1780 1557 1820 1563
rect 2516 1557 2556 1563
rect -19 1537 -13 1543
rect 324 1537 428 1543
rect 436 1537 524 1543
rect 740 1537 876 1543
rect 884 1537 1100 1543
rect 1108 1537 1164 1543
rect 1172 1537 1196 1543
rect 1732 1537 1772 1543
rect 1844 1537 1932 1543
rect 2452 1537 2508 1543
rect 52 1517 92 1523
rect 100 1517 204 1523
rect 212 1517 444 1523
rect 548 1517 780 1523
rect 932 1517 1068 1523
rect 1076 1517 1132 1523
rect 1252 1517 1740 1523
rect 1924 1517 1964 1523
rect 1972 1517 1996 1523
rect 2004 1517 2460 1523
rect -19 1497 140 1503
rect 180 1497 204 1503
rect 244 1497 284 1503
rect 292 1497 348 1503
rect 772 1497 956 1503
rect 964 1497 1148 1503
rect 1156 1497 1324 1503
rect 1380 1497 1436 1503
rect 1780 1497 1932 1503
rect 2468 1497 2524 1503
rect 260 1477 284 1483
rect 292 1477 300 1483
rect 756 1477 924 1483
rect 1092 1477 1292 1483
rect 1908 1477 2284 1483
rect 2404 1477 2652 1483
rect -19 1457 12 1463
rect 84 1457 108 1463
rect 116 1457 316 1463
rect 468 1457 604 1463
rect 612 1457 636 1463
rect 820 1457 1004 1463
rect 1012 1457 1084 1463
rect 1124 1457 1228 1463
rect 1924 1457 2252 1463
rect 2260 1457 2732 1463
rect 212 1437 700 1443
rect 900 1437 1068 1443
rect 1540 1417 1580 1423
rect 2072 1414 2120 1416
rect 2072 1406 2076 1414
rect 2086 1406 2092 1414
rect 2100 1406 2106 1414
rect 2116 1406 2120 1414
rect 2072 1404 2120 1406
rect 324 1397 444 1403
rect 452 1397 556 1403
rect 564 1397 652 1403
rect 1396 1397 1484 1403
rect 2596 1397 2636 1403
rect 2740 1397 2780 1403
rect 308 1377 476 1383
rect 1860 1377 2044 1383
rect 2052 1377 2076 1383
rect 180 1357 268 1363
rect 372 1357 556 1363
rect 580 1357 716 1363
rect 756 1357 780 1363
rect 1460 1357 1564 1363
rect 1732 1357 1996 1363
rect 2004 1357 2220 1363
rect 2292 1357 2412 1363
rect 2484 1357 2540 1363
rect 388 1337 460 1343
rect 468 1337 492 1343
rect 1028 1337 1068 1343
rect 1076 1337 1116 1343
rect 1700 1337 1884 1343
rect 1892 1337 2124 1343
rect 2164 1337 2204 1343
rect 2468 1337 2812 1343
rect 52 1317 108 1323
rect 516 1317 620 1323
rect 836 1317 1228 1323
rect 1236 1317 1372 1323
rect 1780 1317 1820 1323
rect 1956 1317 2028 1323
rect 2436 1317 2540 1323
rect 2564 1317 2588 1323
rect 2660 1317 2700 1323
rect -19 1297 12 1303
rect 1060 1297 1132 1303
rect 1140 1297 1196 1303
rect 1204 1297 1244 1303
rect 1284 1297 1628 1303
rect 1732 1297 2140 1303
rect 2196 1297 2252 1303
rect 2260 1297 2300 1303
rect 2340 1297 2476 1303
rect 2484 1297 2620 1303
rect 724 1277 1084 1283
rect 1156 1277 1212 1283
rect 1828 1277 1836 1283
rect 1844 1277 1852 1283
rect 2388 1277 2508 1283
rect 2973 1277 2979 1283
rect 1796 1257 2348 1263
rect 2468 1257 2492 1263
rect 1572 1237 1596 1243
rect 1700 1217 1884 1223
rect 1892 1217 1980 1223
rect 824 1214 872 1216
rect 824 1206 828 1214
rect 838 1206 844 1214
rect 852 1206 858 1214
rect 868 1206 872 1214
rect 824 1204 872 1206
rect 148 1197 556 1203
rect 2973 1197 2979 1203
rect 308 1177 332 1183
rect 1492 1177 1516 1183
rect 1524 1177 1948 1183
rect 1956 1177 1964 1183
rect 1972 1177 2012 1183
rect 1252 1157 1372 1163
rect 916 1137 1292 1143
rect 1300 1137 1308 1143
rect 1636 1137 2236 1143
rect 2532 1137 2636 1143
rect 692 1117 764 1123
rect 772 1117 812 1123
rect 964 1117 1020 1123
rect 1172 1117 1196 1123
rect 1236 1117 1420 1123
rect 1940 1117 2428 1123
rect 2436 1117 2460 1123
rect 2500 1117 2556 1123
rect 2580 1117 2604 1123
rect 260 1097 380 1103
rect 804 1097 988 1103
rect 996 1097 1036 1103
rect 1044 1097 1052 1103
rect 1060 1097 1260 1103
rect 1268 1097 1356 1103
rect 2148 1097 2172 1103
rect 2404 1097 2444 1103
rect 2477 1097 2508 1103
rect 500 1077 700 1083
rect 1156 1077 1180 1083
rect 1188 1077 1228 1083
rect 1236 1077 1260 1083
rect 1332 1077 1452 1083
rect 1716 1077 1740 1083
rect 1748 1077 1804 1083
rect 2180 1077 2284 1083
rect 2292 1077 2300 1083
rect 2477 1083 2483 1097
rect 2516 1097 2588 1103
rect 2436 1077 2483 1083
rect 2500 1077 2780 1083
rect 1076 1057 1324 1063
rect 1364 1057 1724 1063
rect 2164 1057 2220 1063
rect 2276 1057 2668 1063
rect 532 1037 764 1043
rect 1396 1037 1580 1043
rect 1988 1037 2428 1043
rect 2436 1037 2476 1043
rect 2484 1037 2524 1043
rect 500 1017 812 1023
rect 820 1017 1068 1023
rect 1124 1017 1436 1023
rect 1444 1017 1484 1023
rect 1492 1017 1532 1023
rect 2340 1017 2348 1023
rect 2072 1014 2120 1016
rect 2072 1006 2076 1014
rect 2086 1006 2092 1014
rect 2100 1006 2106 1014
rect 2116 1006 2120 1014
rect 2072 1004 2120 1006
rect 564 997 716 1003
rect 1108 977 1196 983
rect 2036 977 2044 983
rect 2973 977 2979 983
rect 372 957 460 963
rect 468 957 556 963
rect 1636 957 1884 963
rect 1924 957 1980 963
rect 2036 957 2140 963
rect 2148 957 2188 963
rect 2196 957 2412 963
rect 2468 957 2508 963
rect 148 937 348 943
rect 740 937 1084 943
rect 1652 937 1788 943
rect 1972 937 2284 943
rect 2484 937 2796 943
rect 452 917 1036 923
rect 1044 917 1068 923
rect 1492 917 1532 923
rect 1828 917 1916 923
rect 2036 917 2172 923
rect 2276 917 2492 923
rect 852 897 1180 903
rect 1556 897 1676 903
rect 1876 897 1916 903
rect 2052 897 2236 903
rect 2244 897 2268 903
rect 2276 897 2300 903
rect 2324 897 2444 903
rect 2452 897 2604 903
rect 436 877 476 883
rect 484 877 524 883
rect 532 877 1100 883
rect 1108 877 1132 883
rect 1252 877 1276 883
rect 1604 877 1660 883
rect 1716 877 1740 883
rect 1748 877 1772 883
rect 1780 877 1804 883
rect 1812 877 2092 883
rect 2100 877 2156 883
rect 2372 877 2412 883
rect 2420 877 2476 883
rect 2484 877 2556 883
rect 340 857 412 863
rect 420 857 988 863
rect 1588 857 1804 863
rect 1812 857 1932 863
rect 1940 857 2220 863
rect 2436 857 2460 863
rect -19 837 -13 843
rect 2196 837 2524 843
rect 2532 837 2620 843
rect 708 817 764 823
rect 824 814 872 816
rect 824 806 828 814
rect 838 806 844 814
rect 852 806 858 814
rect 868 806 872 814
rect 824 804 872 806
rect 1556 797 1644 803
rect 596 777 1164 783
rect 1172 777 1452 783
rect 1620 757 2780 763
rect 1012 737 1228 743
rect 1956 737 2156 743
rect 2212 737 2316 743
rect 340 717 412 723
rect 420 717 1276 723
rect 1332 717 1372 723
rect 1380 717 1436 723
rect 1828 717 1852 723
rect 2020 717 2147 723
rect 2141 704 2147 717
rect 2164 717 2428 723
rect 676 697 876 703
rect 980 697 1036 703
rect 1076 697 1116 703
rect 1124 697 1340 703
rect 1860 697 1916 703
rect 1988 697 2028 703
rect 2148 697 2204 703
rect 2436 697 2524 703
rect 148 677 348 683
rect 468 677 508 683
rect 516 677 572 683
rect 868 677 1020 683
rect 1092 677 1132 683
rect 1300 677 1788 683
rect 1828 677 1916 683
rect 2004 677 2044 683
rect 2052 677 2092 683
rect 2564 677 2812 683
rect 1133 664 1139 676
rect 180 657 508 663
rect 516 657 700 663
rect 1140 657 1324 663
rect 1892 657 2348 663
rect 2068 637 2140 643
rect 2372 617 2828 623
rect 2072 614 2120 616
rect 2072 606 2076 614
rect 2086 606 2092 614
rect 2100 606 2106 614
rect 2116 606 2120 614
rect 2072 604 2120 606
rect 500 577 748 583
rect 788 577 924 583
rect 1780 577 1836 583
rect 1844 577 1916 583
rect 1924 577 2236 583
rect 2244 577 2300 583
rect 2308 577 2588 583
rect 2596 577 2636 583
rect 2852 577 2876 583
rect 596 557 684 563
rect 724 557 1052 563
rect 1396 557 1644 563
rect 2004 557 2188 563
rect 2292 557 2332 563
rect 2884 557 2924 563
rect 2973 557 2979 563
rect 148 537 348 543
rect 564 537 620 543
rect 628 537 828 543
rect 1156 537 1308 543
rect 1364 537 1420 543
rect 1428 537 1612 543
rect 1908 537 2156 543
rect 2324 537 2412 543
rect 2436 537 2460 543
rect 2468 537 2556 543
rect 2660 537 2748 543
rect 2756 537 2828 543
rect 2836 537 2892 543
rect 452 517 588 523
rect 644 517 700 523
rect 772 517 1260 523
rect 1380 517 1452 523
rect 1748 517 1788 523
rect 1796 517 1852 523
rect 2020 517 2028 523
rect 2196 517 2364 523
rect 2372 517 2524 523
rect 2564 517 2604 523
rect 2612 517 2668 523
rect 2724 517 2764 523
rect 372 497 652 503
rect 660 497 732 503
rect 740 497 908 503
rect 1172 497 1884 503
rect 2013 503 2019 516
rect 1892 497 2396 503
rect 2404 497 2780 503
rect 2788 497 2892 503
rect 436 477 476 483
rect 1732 477 1868 483
rect 1876 477 1996 483
rect 2484 477 2796 483
rect 2804 477 2908 483
rect 340 457 396 463
rect 1252 457 1356 463
rect 1364 457 1836 463
rect 1892 457 1916 463
rect 1972 457 2268 463
rect 2580 457 2716 463
rect 1956 437 2204 443
rect 2420 437 2476 443
rect 2516 437 2652 443
rect 1588 417 1932 423
rect 2388 417 2700 423
rect 824 414 872 416
rect 824 406 828 414
rect 838 406 844 414
rect 852 406 858 414
rect 868 406 872 414
rect 824 404 872 406
rect 1940 397 2124 403
rect 2484 397 2588 403
rect 868 377 940 383
rect 2084 377 2124 383
rect 2244 377 2508 383
rect 2548 377 2780 383
rect 884 357 1020 363
rect 2308 357 2428 363
rect 2516 357 2652 363
rect 2260 337 2364 343
rect 2372 337 2492 343
rect 340 317 412 323
rect 420 317 508 323
rect 948 317 1068 323
rect 1076 317 1132 323
rect 2164 317 2444 323
rect 2500 317 2556 323
rect 2564 317 2860 323
rect 260 297 636 303
rect 1028 297 1052 303
rect 1700 297 1852 303
rect 2260 297 2300 303
rect 2500 297 2572 303
rect 148 277 348 283
rect 756 277 956 283
rect 1124 277 1132 283
rect 1140 277 1164 283
rect 1316 277 1740 283
rect 2308 277 2364 283
rect 2372 277 2588 283
rect 2740 277 2860 283
rect 612 257 652 263
rect 1309 263 1315 276
rect 660 257 1315 263
rect 1620 257 1852 263
rect 1860 257 1964 263
rect 1972 257 2044 263
rect 2212 257 2316 263
rect 2324 257 2380 263
rect 2468 257 2764 263
rect 180 237 540 243
rect 548 237 780 243
rect 788 237 876 243
rect 2692 217 2764 223
rect 2072 214 2120 216
rect 2072 206 2076 214
rect 2086 206 2092 214
rect 2100 206 2106 214
rect 2116 206 2120 214
rect 2072 204 2120 206
rect 868 197 956 203
rect 1268 197 1292 203
rect 1572 197 1612 203
rect 2500 197 2540 203
rect 2596 197 2636 203
rect -19 177 -13 183
rect 1076 177 1148 183
rect 1156 177 1388 183
rect 2228 177 2716 183
rect 2724 177 2812 183
rect 452 157 492 163
rect 1172 157 1276 163
rect 2052 157 2460 163
rect 2644 157 2764 163
rect 148 137 348 143
rect 404 137 444 143
rect 468 137 508 143
rect 852 137 1052 143
rect 1108 137 1180 143
rect 1188 137 1292 143
rect 1396 137 1596 143
rect 2020 137 2284 143
rect 2612 137 2636 143
rect 2644 137 2732 143
rect 340 117 444 123
rect 1108 117 1196 123
rect 2132 117 2380 123
rect 2628 117 2684 123
rect 2836 117 2940 123
rect -19 97 -13 103
rect 1044 97 1212 103
rect 1284 97 1324 103
rect 1332 97 1404 103
rect 2548 97 2668 103
rect 2676 97 2780 103
rect 2868 97 2892 103
rect 2388 77 2764 83
rect 824 14 872 16
rect 824 6 828 14
rect 838 6 844 14
rect 852 6 858 14
rect 868 6 872 14
rect 824 4 872 6
<< m4contact >>
rect 828 2006 830 2014
rect 830 2006 836 2014
rect 844 2006 852 2014
rect 860 2006 866 2014
rect 866 2006 868 2014
rect 108 1896 116 1904
rect 300 1896 308 1904
rect 1132 1876 1140 1884
rect 300 1856 308 1864
rect 2508 1856 2516 1864
rect 780 1816 788 1824
rect 2076 1806 2078 1814
rect 2078 1806 2084 1814
rect 2092 1806 2100 1814
rect 2108 1806 2114 1814
rect 2114 1806 2116 1814
rect 2380 1736 2388 1744
rect 2380 1696 2388 1704
rect 1132 1636 1140 1644
rect 828 1606 830 1614
rect 830 1606 836 1614
rect 844 1606 852 1614
rect 860 1606 866 1614
rect 866 1606 868 1614
rect 300 1476 308 1484
rect 2764 1476 2772 1484
rect 108 1456 116 1464
rect 2076 1406 2078 1414
rect 2078 1406 2084 1414
rect 2092 1406 2100 1414
rect 2108 1406 2114 1414
rect 2114 1406 2116 1414
rect 1484 1396 1492 1404
rect 2636 1396 2644 1404
rect 780 1356 788 1364
rect 2540 1356 2548 1364
rect 460 1336 468 1344
rect 2348 1256 2356 1264
rect 828 1206 830 1214
rect 830 1206 836 1214
rect 844 1206 852 1214
rect 860 1206 866 1214
rect 866 1206 868 1214
rect 300 1176 308 1184
rect 1484 1176 1492 1184
rect 2604 1116 2612 1124
rect 1740 1076 1748 1084
rect 2348 1016 2356 1024
rect 2076 1006 2078 1014
rect 2078 1006 2084 1014
rect 2092 1006 2100 1014
rect 2108 1006 2114 1014
rect 2114 1006 2116 1014
rect 2028 976 2036 984
rect 460 956 468 964
rect 828 806 830 814
rect 830 806 836 814
rect 844 806 852 814
rect 860 806 866 814
rect 866 806 868 814
rect 1132 656 1140 664
rect 2076 606 2078 614
rect 2078 606 2084 614
rect 2092 606 2100 614
rect 2108 606 2114 614
rect 2114 606 2116 614
rect 2028 516 2036 524
rect 1164 496 1172 504
rect 828 406 830 414
rect 830 406 836 414
rect 844 406 852 414
rect 860 406 866 414
rect 866 406 868 414
rect 2508 356 2516 364
rect 1164 296 1172 304
rect 1132 276 1140 284
rect 1740 276 1748 284
rect 2764 216 2772 224
rect 2076 206 2078 214
rect 2078 206 2084 214
rect 2092 206 2100 214
rect 2108 206 2114 214
rect 2114 206 2116 214
rect 2636 156 2644 164
rect 1740 136 1748 144
rect 2604 136 2612 144
rect 2540 96 2548 104
rect 2380 76 2388 84
rect 828 6 830 14
rect 830 6 836 14
rect 844 6 852 14
rect 860 6 866 14
rect 866 6 868 14
<< metal4 >>
rect 824 2014 872 2040
rect 824 2006 828 2014
rect 836 2006 844 2014
rect 852 2006 860 2014
rect 868 2006 872 2014
rect 106 1904 118 1906
rect 106 1896 108 1904
rect 116 1896 118 1904
rect 106 1464 118 1896
rect 106 1456 108 1464
rect 116 1456 118 1464
rect 106 1454 118 1456
rect 298 1904 310 1906
rect 298 1896 300 1904
rect 308 1896 310 1904
rect 298 1864 310 1896
rect 298 1856 300 1864
rect 308 1856 310 1864
rect 298 1484 310 1856
rect 298 1476 300 1484
rect 308 1476 310 1484
rect 298 1184 310 1476
rect 778 1824 790 1826
rect 778 1816 780 1824
rect 788 1816 790 1824
rect 778 1364 790 1816
rect 778 1356 780 1364
rect 788 1356 790 1364
rect 778 1354 790 1356
rect 824 1614 872 2006
rect 1130 1884 1142 1886
rect 1130 1876 1132 1884
rect 1140 1876 1142 1884
rect 1130 1644 1142 1876
rect 1130 1636 1132 1644
rect 1140 1636 1142 1644
rect 1130 1634 1142 1636
rect 2072 1814 2120 2040
rect 2072 1806 2076 1814
rect 2084 1806 2092 1814
rect 2100 1806 2108 1814
rect 2116 1806 2120 1814
rect 824 1606 828 1614
rect 836 1606 844 1614
rect 852 1606 860 1614
rect 868 1606 872 1614
rect 298 1176 300 1184
rect 308 1176 310 1184
rect 298 1174 310 1176
rect 458 1344 470 1346
rect 458 1336 460 1344
rect 468 1336 470 1344
rect 458 964 470 1336
rect 458 956 460 964
rect 468 956 470 964
rect 458 954 470 956
rect 824 1214 872 1606
rect 2072 1414 2120 1806
rect 2506 1864 2518 1866
rect 2506 1856 2508 1864
rect 2516 1856 2518 1864
rect 2072 1406 2076 1414
rect 2084 1406 2092 1414
rect 2100 1406 2108 1414
rect 2116 1406 2120 1414
rect 824 1206 828 1214
rect 836 1206 844 1214
rect 852 1206 860 1214
rect 868 1206 872 1214
rect 824 814 872 1206
rect 1482 1404 1494 1406
rect 1482 1396 1484 1404
rect 1492 1396 1494 1404
rect 1482 1184 1494 1396
rect 1482 1176 1484 1184
rect 1492 1176 1494 1184
rect 1482 1174 1494 1176
rect 824 806 828 814
rect 836 806 844 814
rect 852 806 860 814
rect 868 806 872 814
rect 824 414 872 806
rect 1738 1084 1750 1086
rect 1738 1076 1740 1084
rect 1748 1076 1750 1084
rect 824 406 828 414
rect 836 406 844 414
rect 852 406 860 414
rect 868 406 872 414
rect 824 14 872 406
rect 1130 664 1142 666
rect 1130 656 1132 664
rect 1140 656 1142 664
rect 1130 284 1142 656
rect 1162 504 1174 506
rect 1162 496 1164 504
rect 1172 496 1174 504
rect 1162 304 1174 496
rect 1162 296 1164 304
rect 1172 296 1174 304
rect 1162 294 1174 296
rect 1130 276 1132 284
rect 1140 276 1142 284
rect 1130 274 1142 276
rect 1738 284 1750 1076
rect 2072 1014 2120 1406
rect 2378 1744 2390 1746
rect 2378 1736 2380 1744
rect 2388 1736 2390 1744
rect 2378 1704 2390 1736
rect 2378 1696 2380 1704
rect 2388 1696 2390 1704
rect 2346 1264 2358 1266
rect 2346 1256 2348 1264
rect 2356 1256 2358 1264
rect 2346 1024 2358 1256
rect 2346 1016 2348 1024
rect 2356 1016 2358 1024
rect 2346 1014 2358 1016
rect 2072 1006 2076 1014
rect 2084 1006 2092 1014
rect 2100 1006 2108 1014
rect 2116 1006 2120 1014
rect 2026 984 2038 986
rect 2026 976 2028 984
rect 2036 976 2038 984
rect 2026 524 2038 976
rect 2026 516 2028 524
rect 2036 516 2038 524
rect 2026 514 2038 516
rect 2072 614 2120 1006
rect 2072 606 2076 614
rect 2084 606 2092 614
rect 2100 606 2108 614
rect 2116 606 2120 614
rect 1738 276 1740 284
rect 1748 276 1750 284
rect 1738 144 1750 276
rect 1738 136 1740 144
rect 1748 136 1750 144
rect 1738 134 1750 136
rect 2072 214 2120 606
rect 2072 206 2076 214
rect 2084 206 2092 214
rect 2100 206 2108 214
rect 2116 206 2120 214
rect 824 6 828 14
rect 836 6 844 14
rect 852 6 860 14
rect 868 6 872 14
rect 824 -40 872 6
rect 2072 -40 2120 206
rect 2378 84 2390 1696
rect 2506 364 2518 1856
rect 2762 1484 2774 1486
rect 2762 1476 2764 1484
rect 2772 1476 2774 1484
rect 2634 1404 2646 1406
rect 2634 1396 2636 1404
rect 2644 1396 2646 1404
rect 2506 356 2508 364
rect 2516 356 2518 364
rect 2506 354 2518 356
rect 2538 1364 2550 1366
rect 2538 1356 2540 1364
rect 2548 1356 2550 1364
rect 2538 104 2550 1356
rect 2602 1124 2614 1126
rect 2602 1116 2604 1124
rect 2612 1116 2614 1124
rect 2602 144 2614 1116
rect 2634 164 2646 1396
rect 2762 224 2774 1476
rect 2762 216 2764 224
rect 2772 216 2774 224
rect 2762 214 2774 216
rect 2634 156 2636 164
rect 2644 156 2646 164
rect 2634 154 2646 156
rect 2602 136 2604 144
rect 2612 136 2614 144
rect 2602 134 2614 136
rect 2538 96 2540 104
rect 2548 96 2550 104
rect 2538 94 2550 96
rect 2378 76 2380 84
rect 2388 76 2390 84
rect 2378 74 2390 76
use INVX1  INVX1_20
timestamp 1744796300
transform 1 0 8 0 1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_55
timestamp 1744796300
transform 1 0 40 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_39
timestamp 1744796300
transform 1 0 104 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_46
timestamp 1744796300
transform 1 0 152 0 1 1810
box -4 -6 68 206
use NOR2X1  NOR2X1_40
timestamp 1744796300
transform -1 0 264 0 1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_25
timestamp 1744796300
transform 1 0 264 0 1 1810
box -4 -6 68 206
use INVX1  INVX1_21
timestamp 1744796300
transform -1 0 360 0 1 1810
box -4 -6 36 206
use BUFX2  BUFX2_6
timestamp 1744796300
transform 1 0 360 0 1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_25
timestamp 1744796300
transform -1 0 456 0 1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_57
timestamp 1744796300
transform -1 0 520 0 1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_48
timestamp 1744796300
transform 1 0 520 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_26
timestamp 1744796300
transform -1 0 632 0 1 1810
box -4 -6 52 206
use BUFX2  BUFX2_7
timestamp 1744796300
transform 1 0 632 0 1 1810
box -4 -6 52 206
use FILL  FILL_9_0_0
timestamp 1744796300
transform -1 0 696 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_1
timestamp 1744796300
transform -1 0 712 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_0_2
timestamp 1744796300
transform -1 0 728 0 1 1810
box -4 -6 20 206
use DFFSR  DFFSR_3
timestamp 1744796300
transform -1 0 1080 0 1 1810
box -4 -6 356 206
use AOI22X1  AOI22X1_1
timestamp 1744796300
transform 1 0 1080 0 1 1810
box -4 -6 84 206
use INVX1  INVX1_14
timestamp 1744796300
transform -1 0 1192 0 1 1810
box -4 -6 36 206
use BUFX2  BUFX2_3
timestamp 1744796300
transform 1 0 1192 0 1 1810
box -4 -6 52 206
use DFFSR  DFFSR_4
timestamp 1744796300
transform -1 0 1592 0 1 1810
box -4 -6 356 206
use DFFSR  DFFSR_13
timestamp 1744796300
transform 1 0 1592 0 1 1810
box -4 -6 356 206
use FILL  FILL_9_1_0
timestamp 1744796300
transform -1 0 1960 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_1
timestamp 1744796300
transform -1 0 1976 0 1 1810
box -4 -6 20 206
use FILL  FILL_9_1_2
timestamp 1744796300
transform -1 0 1992 0 1 1810
box -4 -6 20 206
use DFFSR  DFFSR_11
timestamp 1744796300
transform -1 0 2344 0 1 1810
box -4 -6 356 206
use OR2X2  OR2X2_1
timestamp 1744796300
transform -1 0 2408 0 1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_10
timestamp 1744796300
transform -1 0 2456 0 1 1810
box -4 -6 52 206
use XOR2X1  XOR2X1_1
timestamp 1744796300
transform 1 0 2456 0 1 1810
box -4 -6 116 206
use DFFSR  DFFSR_9
timestamp 1744796300
transform -1 0 2920 0 1 1810
box -4 -6 356 206
use FILL  FILL_10_1
timestamp 1744796300
transform 1 0 2920 0 1 1810
box -4 -6 20 206
use FILL  FILL_10_2
timestamp 1744796300
transform 1 0 2936 0 1 1810
box -4 -6 20 206
use INVX1  INVX1_17
timestamp 1744796300
transform 1 0 8 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_56
timestamp 1744796300
transform -1 0 104 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_22
timestamp 1744796300
transform -1 0 136 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_53
timestamp 1744796300
transform -1 0 200 0 -1 1810
box -4 -6 68 206
use NAND2X1  NAND2X1_24
timestamp 1744796300
transform 1 0 200 0 -1 1810
box -4 -6 52 206
use OAI21X1  OAI21X1_50
timestamp 1744796300
transform -1 0 312 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_47
timestamp 1744796300
transform -1 0 376 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_52
timestamp 1744796300
transform -1 0 440 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_16
timestamp 1744796300
transform -1 0 472 0 -1 1810
box -4 -6 36 206
use NOR2X1  NOR2X1_41
timestamp 1744796300
transform -1 0 520 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_27
timestamp 1744796300
transform -1 0 568 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_38
timestamp 1744796300
transform 1 0 568 0 -1 1810
box -4 -6 52 206
use NAND2X1  NAND2X1_22
timestamp 1744796300
transform 1 0 616 0 -1 1810
box -4 -6 52 206
use NOR2X1  NOR2X1_37
timestamp 1744796300
transform -1 0 712 0 -1 1810
box -4 -6 52 206
use INVX1  INVX1_1
timestamp 1744796300
transform 1 0 712 0 -1 1810
box -4 -6 36 206
use OR2X2  OR2X2_3
timestamp 1744796300
transform 1 0 744 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_0_0
timestamp 1744796300
transform 1 0 808 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_1
timestamp 1744796300
transform 1 0 824 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_0_2
timestamp 1744796300
transform 1 0 840 0 -1 1810
box -4 -6 20 206
use OAI21X1  OAI21X1_58
timestamp 1744796300
transform 1 0 856 0 -1 1810
box -4 -6 68 206
use OAI21X1  OAI21X1_59
timestamp 1744796300
transform -1 0 984 0 -1 1810
box -4 -6 68 206
use DFFSR  DFFSR_7
timestamp 1744796300
transform -1 0 1336 0 -1 1810
box -4 -6 356 206
use DFFSR  DFFSR_12
timestamp 1744796300
transform 1 0 1336 0 -1 1810
box -4 -6 356 206
use OAI21X1  OAI21X1_8
timestamp 1744796300
transform -1 0 1752 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_8
timestamp 1744796300
transform 1 0 1752 0 -1 1810
box -4 -6 36 206
use NAND2X1  NAND2X1_11
timestamp 1744796300
transform -1 0 1832 0 -1 1810
box -4 -6 52 206
use NAND3X1  NAND3X1_7
timestamp 1744796300
transform 1 0 1832 0 -1 1810
box -4 -6 68 206
use INVX1  INVX1_7
timestamp 1744796300
transform 1 0 1896 0 -1 1810
box -4 -6 36 206
use NAND3X1  NAND3X1_5
timestamp 1744796300
transform -1 0 1992 0 -1 1810
box -4 -6 68 206
use INVX2  INVX2_4
timestamp 1744796300
transform 1 0 1992 0 -1 1810
box -4 -6 36 206
use OAI21X1  OAI21X1_7
timestamp 1744796300
transform -1 0 2088 0 -1 1810
box -4 -6 68 206
use FILL  FILL_8_1_0
timestamp 1744796300
transform 1 0 2088 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_1
timestamp 1744796300
transform 1 0 2104 0 -1 1810
box -4 -6 20 206
use FILL  FILL_8_1_2
timestamp 1744796300
transform 1 0 2120 0 -1 1810
box -4 -6 20 206
use NOR3X1  NOR3X1_1
timestamp 1744796300
transform 1 0 2136 0 -1 1810
box -4 -6 132 206
use OAI21X1  OAI21X1_6
timestamp 1744796300
transform -1 0 2328 0 -1 1810
box -4 -6 68 206
use XNOR2X1  XNOR2X1_1
timestamp 1744796300
transform -1 0 2440 0 -1 1810
box -4 -6 116 206
use OAI21X1  OAI21X1_4
timestamp 1744796300
transform 1 0 2440 0 -1 1810
box -4 -6 68 206
use NAND3X1  NAND3X1_4
timestamp 1744796300
transform -1 0 2568 0 -1 1810
box -4 -6 68 206
use DFFSR  DFFSR_10
timestamp 1744796300
transform -1 0 2920 0 -1 1810
box -4 -6 356 206
use FILL  FILL_9_1
timestamp 1744796300
transform -1 0 2936 0 -1 1810
box -4 -6 20 206
use FILL  FILL_9_2
timestamp 1744796300
transform -1 0 2952 0 -1 1810
box -4 -6 20 206
use INVX1  INVX1_15
timestamp 1744796300
transform 1 0 8 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_28
timestamp 1744796300
transform 1 0 40 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_54
timestamp 1744796300
transform -1 0 152 0 1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_51
timestamp 1744796300
transform 1 0 152 0 1 1410
box -4 -6 68 206
use INVX1  INVX1_19
timestamp 1744796300
transform -1 0 248 0 1 1410
box -4 -6 36 206
use INVX2  INVX2_9
timestamp 1744796300
transform 1 0 248 0 1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_1
timestamp 1744796300
transform 1 0 280 0 1 1410
box -4 -6 52 206
use AOI21X1  AOI21X1_6
timestamp 1744796300
transform 1 0 328 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_1
timestamp 1744796300
transform 1 0 392 0 1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_49
timestamp 1744796300
transform 1 0 440 0 1 1410
box -4 -6 68 206
use NOR2X1  NOR2X1_42
timestamp 1744796300
transform -1 0 552 0 1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_23
timestamp 1744796300
transform 1 0 552 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_43
timestamp 1744796300
transform -1 0 648 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_18
timestamp 1744796300
transform 1 0 648 0 1 1410
box -4 -6 36 206
use AOI22X1  AOI22X1_2
timestamp 1744796300
transform -1 0 760 0 1 1410
box -4 -6 84 206
use OAI21X1  OAI21X1_45
timestamp 1744796300
transform -1 0 824 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_0_0
timestamp 1744796300
transform -1 0 840 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_1
timestamp 1744796300
transform -1 0 856 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_0_2
timestamp 1744796300
transform -1 0 872 0 1 1410
box -4 -6 20 206
use NAND2X1  NAND2X1_20
timestamp 1744796300
transform -1 0 920 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_2
timestamp 1744796300
transform 1 0 920 0 1 1410
box -4 -6 36 206
use NAND2X1  NAND2X1_2
timestamp 1744796300
transform 1 0 952 0 1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_36
timestamp 1744796300
transform 1 0 1000 0 1 1410
box -4 -6 52 206
use OAI22X1  OAI22X1_2
timestamp 1744796300
transform -1 0 1128 0 1 1410
box -4 -6 84 206
use NAND3X1  NAND3X1_24
timestamp 1744796300
transform 1 0 1128 0 1 1410
box -4 -6 68 206
use INVX2  INVX2_8
timestamp 1744796300
transform -1 0 1224 0 1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_43
timestamp 1744796300
transform 1 0 1224 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_21
timestamp 1744796300
transform -1 0 1336 0 1 1410
box -4 -6 52 206
use BUFX4  BUFX4_11
timestamp 1744796300
transform -1 0 1400 0 1 1410
box -4 -6 68 206
use DFFSR  DFFSR_18
timestamp 1744796300
transform 1 0 1400 0 1 1410
box -4 -6 356 206
use OAI21X1  OAI21X1_9
timestamp 1744796300
transform 1 0 1752 0 1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_13
timestamp 1744796300
transform -1 0 1864 0 1 1410
box -4 -6 52 206
use INVX1  INVX1_9
timestamp 1744796300
transform -1 0 1896 0 1 1410
box -4 -6 36 206
use NAND3X1  NAND3X1_8
timestamp 1744796300
transform 1 0 1896 0 1 1410
box -4 -6 68 206
use BUFX4  BUFX4_13
timestamp 1744796300
transform 1 0 1960 0 1 1410
box -4 -6 68 206
use FILL  FILL_7_1_0
timestamp 1744796300
transform -1 0 2040 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_1
timestamp 1744796300
transform -1 0 2056 0 1 1410
box -4 -6 20 206
use FILL  FILL_7_1_2
timestamp 1744796300
transform -1 0 2072 0 1 1410
box -4 -6 20 206
use DFFSR  DFFSR_14
timestamp 1744796300
transform -1 0 2424 0 1 1410
box -4 -6 356 206
use NAND3X1  NAND3X1_3
timestamp 1744796300
transform -1 0 2488 0 1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_1
timestamp 1744796300
transform -1 0 2552 0 1 1410
box -4 -6 68 206
use DFFSR  DFFSR_8
timestamp 1744796300
transform -1 0 2904 0 1 1410
box -4 -6 356 206
use FILL  FILL_8_1
timestamp 1744796300
transform 1 0 2904 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_2
timestamp 1744796300
transform 1 0 2920 0 1 1410
box -4 -6 20 206
use FILL  FILL_8_3
timestamp 1744796300
transform 1 0 2936 0 1 1410
box -4 -6 20 206
use BUFX2  BUFX2_5
timestamp 1744796300
transform -1 0 56 0 -1 1410
box -4 -6 52 206
use INVX2  INVX2_1
timestamp 1744796300
transform 1 0 56 0 -1 1410
box -4 -6 36 206
use DFFSR  DFFSR_1
timestamp 1744796300
transform -1 0 440 0 -1 1410
box -4 -6 356 206
use AOI21X1  AOI21X1_5
timestamp 1744796300
transform 1 0 440 0 -1 1410
box -4 -6 68 206
use AOI22X1  AOI22X1_3
timestamp 1744796300
transform 1 0 504 0 -1 1410
box -4 -6 84 206
use DFFSR  DFFSR_38
timestamp 1744796300
transform 1 0 584 0 -1 1410
box -4 -6 356 206
use FILL  FILL_6_0_0
timestamp 1744796300
transform -1 0 952 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_1
timestamp 1744796300
transform -1 0 968 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_0_2
timestamp 1744796300
transform -1 0 984 0 -1 1410
box -4 -6 20 206
use INVX1  INVX1_3
timestamp 1744796300
transform -1 0 1016 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_35
timestamp 1744796300
transform 1 0 1016 0 -1 1410
box -4 -6 52 206
use NOR2X1  NOR2X1_2
timestamp 1744796300
transform -1 0 1112 0 -1 1410
box -4 -6 52 206
use INVX2  INVX2_7
timestamp 1744796300
transform 1 0 1112 0 -1 1410
box -4 -6 36 206
use OAI21X1  OAI21X1_41
timestamp 1744796300
transform 1 0 1144 0 -1 1410
box -4 -6 68 206
use BUFX4  BUFX4_16
timestamp 1744796300
transform -1 0 1272 0 -1 1410
box -4 -6 68 206
use DFFSR  DFFSR_37
timestamp 1744796300
transform -1 0 1624 0 -1 1410
box -4 -6 356 206
use BUFX4  BUFX4_17
timestamp 1744796300
transform 1 0 1624 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_12
timestamp 1744796300
transform 1 0 1688 0 -1 1410
box -4 -6 52 206
use NAND2X1  NAND2X1_14
timestamp 1744796300
transform 1 0 1736 0 -1 1410
box -4 -6 52 206
use BUFX2  BUFX2_1
timestamp 1744796300
transform 1 0 1784 0 -1 1410
box -4 -6 52 206
use NAND3X1  NAND3X1_9
timestamp 1744796300
transform -1 0 1896 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_10
timestamp 1744796300
transform -1 0 1960 0 -1 1410
box -4 -6 68 206
use XNOR2X1  XNOR2X1_2
timestamp 1744796300
transform 1 0 1960 0 -1 1410
box -4 -6 116 206
use FILL  FILL_6_1_0
timestamp 1744796300
transform 1 0 2072 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_1
timestamp 1744796300
transform 1 0 2088 0 -1 1410
box -4 -6 20 206
use FILL  FILL_6_1_2
timestamp 1744796300
transform 1 0 2104 0 -1 1410
box -4 -6 20 206
use INVX2  INVX2_2
timestamp 1744796300
transform 1 0 2120 0 -1 1410
box -4 -6 36 206
use NOR2X1  NOR2X1_5
timestamp 1744796300
transform -1 0 2200 0 -1 1410
box -4 -6 52 206
use OAI21X1  OAI21X1_11
timestamp 1744796300
transform 1 0 2200 0 -1 1410
box -4 -6 68 206
use NAND2X1  NAND2X1_15
timestamp 1744796300
transform -1 0 2312 0 -1 1410
box -4 -6 52 206
use INVX1  INVX1_6
timestamp 1744796300
transform -1 0 2344 0 -1 1410
box -4 -6 36 206
use BUFX4  BUFX4_2
timestamp 1744796300
transform 1 0 2344 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_12
timestamp 1744796300
transform 1 0 2408 0 -1 1410
box -4 -6 68 206
use NAND3X1  NAND3X1_10
timestamp 1744796300
transform 1 0 2472 0 -1 1410
box -4 -6 68 206
use OAI21X1  OAI21X1_5
timestamp 1744796300
transform 1 0 2536 0 -1 1410
box -4 -6 68 206
use DFFSR  DFFSR_15
timestamp 1744796300
transform -1 0 2952 0 -1 1410
box -4 -6 356 206
use DFFSR  DFFSR_2
timestamp 1744796300
transform 1 0 8 0 1 1010
box -4 -6 356 206
use DFFSR  DFFSR_36
timestamp 1744796300
transform 1 0 360 0 1 1010
box -4 -6 356 206
use NOR2X1  NOR2X1_31
timestamp 1744796300
transform 1 0 712 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_37
timestamp 1744796300
transform -1 0 824 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_0_0
timestamp 1744796300
transform -1 0 840 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_1
timestamp 1744796300
transform -1 0 856 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_0_2
timestamp 1744796300
transform -1 0 872 0 1 1010
box -4 -6 20 206
use NOR2X1  NOR2X1_10
timestamp 1744796300
transform -1 0 920 0 1 1010
box -4 -6 52 206
use NAND2X1  NAND2X1_5
timestamp 1744796300
transform -1 0 968 0 1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_9
timestamp 1744796300
transform -1 0 1016 0 1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_39
timestamp 1744796300
transform -1 0 1080 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_33
timestamp 1744796300
transform -1 0 1128 0 1 1010
box -4 -6 52 206
use BUFX4  BUFX4_6
timestamp 1744796300
transform 1 0 1128 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_42
timestamp 1744796300
transform -1 0 1256 0 1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_38
timestamp 1744796300
transform 1 0 1256 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_3
timestamp 1744796300
transform 1 0 1320 0 1 1010
box -4 -6 52 206
use OAI22X1  OAI22X1_1
timestamp 1744796300
transform -1 0 1448 0 1 1010
box -4 -6 84 206
use NOR2X1  NOR2X1_32
timestamp 1744796300
transform -1 0 1496 0 1 1010
box -4 -6 52 206
use INVX8  INVX8_1
timestamp 1744796300
transform 1 0 1496 0 1 1010
box -4 -6 84 206
use CLKBUF1  CLKBUF1_1
timestamp 1744796300
transform -1 0 1720 0 1 1010
box -4 -6 148 206
use INVX8  INVX8_2
timestamp 1744796300
transform 1 0 1720 0 1 1010
box -4 -6 84 206
use CLKBUF1  CLKBUF1_3
timestamp 1744796300
transform 1 0 1800 0 1 1010
box -4 -6 148 206
use BUFX4  BUFX4_12
timestamp 1744796300
transform 1 0 1944 0 1 1010
box -4 -6 68 206
use BUFX4  BUFX4_14
timestamp 1744796300
transform 1 0 2008 0 1 1010
box -4 -6 68 206
use FILL  FILL_5_1_0
timestamp 1744796300
transform 1 0 2072 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_1
timestamp 1744796300
transform 1 0 2088 0 1 1010
box -4 -6 20 206
use FILL  FILL_5_1_2
timestamp 1744796300
transform 1 0 2104 0 1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_11
timestamp 1744796300
transform 1 0 2120 0 1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_6
timestamp 1744796300
transform -1 0 2232 0 1 1010
box -4 -6 52 206
use BUFX4  BUFX4_19
timestamp 1744796300
transform 1 0 2232 0 1 1010
box -4 -6 68 206
use XNOR2X1  XNOR2X1_3
timestamp 1744796300
transform 1 0 2296 0 1 1010
box -4 -6 116 206
use INVX2  INVX2_3
timestamp 1744796300
transform -1 0 2440 0 1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_13
timestamp 1744796300
transform 1 0 2440 0 1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_12
timestamp 1744796300
transform 1 0 2504 0 1 1010
box -4 -6 68 206
use DFFSR  DFFSR_16
timestamp 1744796300
transform -1 0 2920 0 1 1010
box -4 -6 356 206
use FILL  FILL_6_1
timestamp 1744796300
transform 1 0 2920 0 1 1010
box -4 -6 20 206
use FILL  FILL_6_2
timestamp 1744796300
transform 1 0 2936 0 1 1010
box -4 -6 20 206
use DFFSR  DFFSR_28
timestamp 1744796300
transform 1 0 8 0 -1 1010
box -4 -6 356 206
use NOR2X1  NOR2X1_23
timestamp 1744796300
transform 1 0 360 0 -1 1010
box -4 -6 52 206
use OAI21X1  OAI21X1_29
timestamp 1744796300
transform -1 0 472 0 -1 1010
box -4 -6 68 206
use BUFX4  BUFX4_5
timestamp 1744796300
transform -1 0 536 0 -1 1010
box -4 -6 68 206
use BUFX4  BUFX4_9
timestamp 1744796300
transform -1 0 600 0 -1 1010
box -4 -6 68 206
use DFFSR  DFFSR_39
timestamp 1744796300
transform 1 0 600 0 -1 1010
box -4 -6 356 206
use FILL  FILL_4_0_0
timestamp 1744796300
transform -1 0 968 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_1
timestamp 1744796300
transform -1 0 984 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_0_2
timestamp 1744796300
transform -1 0 1000 0 -1 1010
box -4 -6 20 206
use OAI21X1  OAI21X1_40
timestamp 1744796300
transform -1 0 1064 0 -1 1010
box -4 -6 68 206
use NOR2X1  NOR2X1_34
timestamp 1744796300
transform -1 0 1112 0 -1 1010
box -4 -6 52 206
use BUFX4  BUFX4_7
timestamp 1744796300
transform -1 0 1176 0 -1 1010
box -4 -6 68 206
use DFFSR  DFFSR_6
timestamp 1744796300
transform -1 0 1528 0 -1 1010
box -4 -6 356 206
use OAI21X1  OAI21X1_44
timestamp 1744796300
transform 1 0 1528 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_17
timestamp 1744796300
transform -1 0 1656 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_14
timestamp 1744796300
transform -1 0 1720 0 -1 1010
box -4 -6 68 206
use BUFX2  BUFX2_2
timestamp 1744796300
transform -1 0 1768 0 -1 1010
box -4 -6 52 206
use NOR2X1  NOR2X1_17
timestamp 1744796300
transform 1 0 1768 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_11
timestamp 1744796300
transform 1 0 1816 0 -1 1010
box -4 -6 36 206
use OAI21X1  OAI21X1_16
timestamp 1744796300
transform 1 0 1848 0 -1 1010
box -4 -6 68 206
use INVX1  INVX1_10
timestamp 1744796300
transform 1 0 1912 0 -1 1010
box -4 -6 36 206
use NOR3X1  NOR3X1_2
timestamp 1744796300
transform -1 0 2072 0 -1 1010
box -4 -6 132 206
use FILL  FILL_4_1_0
timestamp 1744796300
transform -1 0 2088 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_1
timestamp 1744796300
transform -1 0 2104 0 -1 1010
box -4 -6 20 206
use FILL  FILL_4_1_2
timestamp 1744796300
transform -1 0 2120 0 -1 1010
box -4 -6 20 206
use NAND3X1  NAND3X1_2
timestamp 1744796300
transform -1 0 2184 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_14
timestamp 1744796300
transform 1 0 2184 0 -1 1010
box -4 -6 68 206
use NAND2X1  NAND2X1_16
timestamp 1744796300
transform 1 0 2248 0 -1 1010
box -4 -6 52 206
use INVX1  INVX1_5
timestamp 1744796300
transform -1 0 2328 0 -1 1010
box -4 -6 36 206
use BUFX4  BUFX4_1
timestamp 1744796300
transform 1 0 2328 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_13
timestamp 1744796300
transform -1 0 2456 0 -1 1010
box -4 -6 68 206
use OAI21X1  OAI21X1_15
timestamp 1744796300
transform -1 0 2520 0 -1 1010
box -4 -6 68 206
use NAND3X1  NAND3X1_17
timestamp 1744796300
transform 1 0 2520 0 -1 1010
box -4 -6 68 206
use DFFSR  DFFSR_17
timestamp 1744796300
transform -1 0 2936 0 -1 1010
box -4 -6 356 206
use FILL  FILL_5_1
timestamp 1744796300
transform -1 0 2952 0 -1 1010
box -4 -6 20 206
use DFFSR  DFFSR_31
timestamp 1744796300
transform 1 0 8 0 1 610
box -4 -6 356 206
use NOR2X1  NOR2X1_26
timestamp 1744796300
transform 1 0 360 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_32
timestamp 1744796300
transform -1 0 472 0 1 610
box -4 -6 68 206
use BUFX4  BUFX4_3
timestamp 1744796300
transform 1 0 472 0 1 610
box -4 -6 68 206
use DFFSR  DFFSR_29
timestamp 1744796300
transform 1 0 536 0 1 610
box -4 -6 356 206
use FILL  FILL_3_0_0
timestamp 1744796300
transform 1 0 888 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_1
timestamp 1744796300
transform 1 0 904 0 1 610
box -4 -6 20 206
use FILL  FILL_3_0_2
timestamp 1744796300
transform 1 0 920 0 1 610
box -4 -6 20 206
use NOR2X1  NOR2X1_24
timestamp 1744796300
transform 1 0 936 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_13
timestamp 1744796300
transform -1 0 1032 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_30
timestamp 1744796300
transform -1 0 1096 0 1 610
box -4 -6 68 206
use BUFX4  BUFX4_4
timestamp 1744796300
transform 1 0 1096 0 1 610
box -4 -6 68 206
use BUFX4  BUFX4_15
timestamp 1744796300
transform -1 0 1224 0 1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_6
timestamp 1744796300
transform -1 0 1272 0 1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_12
timestamp 1744796300
transform 1 0 1272 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_31
timestamp 1744796300
transform 1 0 1320 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_25
timestamp 1744796300
transform -1 0 1432 0 1 610
box -4 -6 52 206
use DFFSR  DFFSR_5
timestamp 1744796300
transform -1 0 1784 0 1 610
box -4 -6 356 206
use NAND2X1  NAND2X1_8
timestamp 1744796300
transform 1 0 1784 0 1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_2
timestamp 1744796300
transform 1 0 1832 0 1 610
box -4 -6 68 206
use INVX2  INVX2_5
timestamp 1744796300
transform -1 0 1928 0 1 610
box -4 -6 36 206
use INVX1  INVX1_4
timestamp 1744796300
transform -1 0 1960 0 1 610
box -4 -6 36 206
use NAND3X1  NAND3X1_16
timestamp 1744796300
transform -1 0 2024 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_2
timestamp 1744796300
transform 1 0 2024 0 1 610
box -4 -6 68 206
use FILL  FILL_3_1_0
timestamp 1744796300
transform 1 0 2088 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_1
timestamp 1744796300
transform 1 0 2104 0 1 610
box -4 -6 20 206
use FILL  FILL_3_1_2
timestamp 1744796300
transform 1 0 2120 0 1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_1
timestamp 1744796300
transform 1 0 2136 0 1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_4
timestamp 1744796300
transform -1 0 2248 0 1 610
box -4 -6 52 206
use AND2X2  AND2X2_1
timestamp 1744796300
transform 1 0 2248 0 1 610
box -4 -6 68 206
use AOI21X1  AOI21X1_1
timestamp 1744796300
transform 1 0 2312 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_19
timestamp 1744796300
transform 1 0 2376 0 1 610
box -4 -6 68 206
use AND2X2  AND2X2_4
timestamp 1744796300
transform 1 0 2440 0 1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_20
timestamp 1744796300
transform 1 0 2504 0 1 610
box -4 -6 68 206
use INVX2  INVX2_6
timestamp 1744796300
transform -1 0 2600 0 1 610
box -4 -6 36 206
use DFFSR  DFFSR_20
timestamp 1744796300
transform -1 0 2952 0 1 610
box -4 -6 356 206
use DFFSR  DFFSR_33
timestamp 1744796300
transform 1 0 8 0 -1 610
box -4 -6 356 206
use NOR2X1  NOR2X1_28
timestamp 1744796300
transform 1 0 360 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_34
timestamp 1744796300
transform -1 0 472 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_4
timestamp 1744796300
transform -1 0 520 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_7
timestamp 1744796300
transform -1 0 568 0 -1 610
box -4 -6 52 206
use OAI21X1  OAI21X1_36
timestamp 1744796300
transform 1 0 568 0 -1 610
box -4 -6 68 206
use BUFX4  BUFX4_8
timestamp 1744796300
transform -1 0 696 0 -1 610
box -4 -6 68 206
use NOR2X1  NOR2X1_30
timestamp 1744796300
transform -1 0 744 0 -1 610
box -4 -6 52 206
use NOR2X1  NOR2X1_11
timestamp 1744796300
transform 1 0 744 0 -1 610
box -4 -6 52 206
use FILL  FILL_2_0_0
timestamp 1744796300
transform -1 0 808 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_1
timestamp 1744796300
transform -1 0 824 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_0_2
timestamp 1744796300
transform -1 0 840 0 -1 610
box -4 -6 20 206
use DFFSR  DFFSR_35
timestamp 1744796300
transform -1 0 1192 0 -1 610
box -4 -6 356 206
use NOR2X1  NOR2X1_16
timestamp 1744796300
transform -1 0 1240 0 -1 610
box -4 -6 52 206
use AND2X2  AND2X2_3
timestamp 1744796300
transform 1 0 1240 0 -1 610
box -4 -6 68 206
use BUFX4  BUFX4_20
timestamp 1744796300
transform -1 0 1368 0 -1 610
box -4 -6 68 206
use BUFX4  BUFX4_10
timestamp 1744796300
transform 1 0 1368 0 -1 610
box -4 -6 68 206
use DFFSR  DFFSR_30
timestamp 1744796300
transform -1 0 1784 0 -1 610
box -4 -6 356 206
use BUFX4  BUFX4_18
timestamp 1744796300
transform -1 0 1848 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_18
timestamp 1744796300
transform -1 0 1912 0 -1 610
box -4 -6 68 206
use OAI21X1  OAI21X1_22
timestamp 1744796300
transform -1 0 1976 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_15
timestamp 1744796300
transform -1 0 2040 0 -1 610
box -4 -6 68 206
use FILL  FILL_2_1_0
timestamp 1744796300
transform -1 0 2056 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_1
timestamp 1744796300
transform -1 0 2072 0 -1 610
box -4 -6 20 206
use FILL  FILL_2_1_2
timestamp 1744796300
transform -1 0 2088 0 -1 610
box -4 -6 20 206
use OAI21X1  OAI21X1_18
timestamp 1744796300
transform -1 0 2152 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_17
timestamp 1744796300
transform -1 0 2200 0 -1 610
box -4 -6 52 206
use OR2X2  OR2X2_2
timestamp 1744796300
transform -1 0 2264 0 -1 610
box -4 -6 68 206
use INVX1  INVX1_13
timestamp 1744796300
transform -1 0 2296 0 -1 610
box -4 -6 36 206
use INVX1  INVX1_12
timestamp 1744796300
transform 1 0 2296 0 -1 610
box -4 -6 36 206
use OAI21X1  OAI21X1_21
timestamp 1744796300
transform -1 0 2392 0 -1 610
box -4 -6 68 206
use NOR3X1  NOR3X1_3
timestamp 1744796300
transform 1 0 2392 0 -1 610
box -4 -6 132 206
use NOR2X1  NOR2X1_19
timestamp 1744796300
transform -1 0 2568 0 -1 610
box -4 -6 52 206
use NAND3X1  NAND3X1_20
timestamp 1744796300
transform 1 0 2568 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_22
timestamp 1744796300
transform 1 0 2632 0 -1 610
box -4 -6 68 206
use AND2X2  AND2X2_2
timestamp 1744796300
transform 1 0 2696 0 -1 610
box -4 -6 68 206
use NAND3X1  NAND3X1_19
timestamp 1744796300
transform 1 0 2760 0 -1 610
box -4 -6 68 206
use NAND2X1  NAND2X1_3
timestamp 1744796300
transform -1 0 2872 0 -1 610
box -4 -6 52 206
use AOI21X1  AOI21X1_4
timestamp 1744796300
transform 1 0 2872 0 -1 610
box -4 -6 68 206
use FILL  FILL_3_1
timestamp 1744796300
transform -1 0 2952 0 -1 610
box -4 -6 20 206
use DFFSR  DFFSR_34
timestamp 1744796300
transform 1 0 8 0 1 210
box -4 -6 356 206
use NOR2X1  NOR2X1_29
timestamp 1744796300
transform 1 0 360 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_35
timestamp 1744796300
transform -1 0 472 0 1 210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_2
timestamp 1744796300
transform -1 0 616 0 1 210
box -4 -6 148 206
use DFFSR  DFFSR_25
timestamp 1744796300
transform 1 0 616 0 1 210
box -4 -6 356 206
use FILL  FILL_1_0_0
timestamp 1744796300
transform -1 0 984 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_1
timestamp 1744796300
transform -1 0 1000 0 1 210
box -4 -6 20 206
use FILL  FILL_1_0_2
timestamp 1744796300
transform -1 0 1016 0 1 210
box -4 -6 20 206
use NOR2X1  NOR2X1_20
timestamp 1744796300
transform -1 0 1064 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_26
timestamp 1744796300
transform -1 0 1128 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_15
timestamp 1744796300
transform 1 0 1128 0 1 210
box -4 -6 52 206
use NAND2X1  NAND2X1_7
timestamp 1744796300
transform -1 0 1224 0 1 210
box -4 -6 52 206
use INVX8  INVX8_3
timestamp 1744796300
transform -1 0 1304 0 1 210
box -4 -6 84 206
use CLKBUF1  CLKBUF1_4
timestamp 1744796300
transform 1 0 1304 0 1 210
box -4 -6 148 206
use DFFSR  DFFSR_21
timestamp 1744796300
transform 1 0 1448 0 1 210
box -4 -6 356 206
use DFFSR  DFFSR_19
timestamp 1744796300
transform 1 0 1800 0 1 210
box -4 -6 356 206
use FILL  FILL_1_1_0
timestamp 1744796300
transform 1 0 2152 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_1
timestamp 1744796300
transform 1 0 2168 0 1 210
box -4 -6 20 206
use FILL  FILL_1_1_2
timestamp 1744796300
transform 1 0 2184 0 1 210
box -4 -6 20 206
use NAND2X1  NAND2X1_19
timestamp 1744796300
transform 1 0 2200 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_24
timestamp 1744796300
transform 1 0 2248 0 1 210
box -4 -6 68 206
use AOI21X1  AOI21X1_3
timestamp 1744796300
transform -1 0 2376 0 1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_21
timestamp 1744796300
transform 1 0 2376 0 1 210
box -4 -6 68 206
use NAND2X1  NAND2X1_18
timestamp 1744796300
transform 1 0 2440 0 1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_23
timestamp 1744796300
transform 1 0 2488 0 1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_18
timestamp 1744796300
transform -1 0 2600 0 1 210
box -4 -6 52 206
use DFFSR  DFFSR_24
timestamp 1744796300
transform 1 0 2600 0 1 210
box -4 -6 356 206
use DFFSR  DFFSR_32
timestamp 1744796300
transform 1 0 8 0 -1 210
box -4 -6 356 206
use NOR2X1  NOR2X1_27
timestamp 1744796300
transform 1 0 360 0 -1 210
box -4 -6 52 206
use NOR2X1  NOR2X1_8
timestamp 1744796300
transform 1 0 408 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_33
timestamp 1744796300
transform -1 0 520 0 -1 210
box -4 -6 68 206
use CLKBUF1  CLKBUF1_5
timestamp 1744796300
transform -1 0 664 0 -1 210
box -4 -6 148 206
use FILL  FILL_0_0_0
timestamp 1744796300
transform 1 0 664 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_1
timestamp 1744796300
transform 1 0 680 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_0_2
timestamp 1744796300
transform 1 0 696 0 -1 210
box -4 -6 20 206
use DFFSR  DFFSR_27
timestamp 1744796300
transform 1 0 712 0 -1 210
box -4 -6 356 206
use NOR2X1  NOR2X1_22
timestamp 1744796300
transform 1 0 1064 0 -1 210
box -4 -6 52 206
use BUFX2  BUFX2_4
timestamp 1744796300
transform -1 0 1160 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_28
timestamp 1744796300
transform 1 0 1160 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_14
timestamp 1744796300
transform 1 0 1224 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_27
timestamp 1744796300
transform 1 0 1272 0 -1 210
box -4 -6 68 206
use NOR2X1  NOR2X1_21
timestamp 1744796300
transform -1 0 1384 0 -1 210
box -4 -6 52 206
use DFFSR  DFFSR_26
timestamp 1744796300
transform -1 0 1736 0 -1 210
box -4 -6 356 206
use CLKBUF1  CLKBUF1_6
timestamp 1744796300
transform 1 0 1736 0 -1 210
box -4 -6 148 206
use DFFSR  DFFSR_23
timestamp 1744796300
transform 1 0 1880 0 -1 210
box -4 -6 356 206
use FILL  FILL_0_1_0
timestamp 1744796300
transform -1 0 2248 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_1
timestamp 1744796300
transform -1 0 2264 0 -1 210
box -4 -6 20 206
use FILL  FILL_0_1_2
timestamp 1744796300
transform -1 0 2280 0 -1 210
box -4 -6 20 206
use DFFSR  DFFSR_22
timestamp 1744796300
transform -1 0 2632 0 -1 210
box -4 -6 356 206
use NAND2X1  NAND2X1_9
timestamp 1744796300
transform 1 0 2632 0 -1 210
box -4 -6 52 206
use OAI21X1  OAI21X1_3
timestamp 1744796300
transform -1 0 2744 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_6
timestamp 1744796300
transform 1 0 2744 0 -1 210
box -4 -6 68 206
use OAI21X1  OAI21X1_25
timestamp 1744796300
transform 1 0 2808 0 -1 210
box -4 -6 68 206
use NAND3X1  NAND3X1_23
timestamp 1744796300
transform 1 0 2872 0 -1 210
box -4 -6 68 206
use FILL  FILL_1_1
timestamp 1744796300
transform -1 0 2952 0 -1 210
box -4 -6 20 206
<< labels >>
flabel metal4 s 824 -40 872 -16 7 FreeSans 24 270 0 0 vdd
port 0 nsew
flabel metal4 s 2072 -40 2120 -16 7 FreeSans 24 270 0 0 gnd
port 1 nsew
flabel metal2 s 1741 -23 1747 -17 7 FreeSans 24 270 0 0 clk
port 2 nsew
flabel metal2 s 1261 -23 1267 -17 7 FreeSans 24 270 0 0 reset
port 3 nsew
flabel metal2 s 605 2037 611 2043 3 FreeSans 24 90 0 0 insert_card
port 4 nsew
flabel metal3 s -19 97 -13 103 7 FreeSans 24 0 0 0 pin_input[0]
port 5 nsew
flabel metal3 s 2973 1197 2979 1203 3 FreeSans 24 0 0 0 pin_input[1]
port 6 nsew
flabel metal2 s 1149 2037 1155 2043 3 FreeSans 24 90 0 0 pin_input[2]
port 7 nsew
flabel metal3 s 2973 1277 2979 1283 3 FreeSans 24 0 0 0 pin_input[3]
port 8 nsew
flabel metal2 s 237 -23 243 -17 7 FreeSans 24 270 0 0 pin_input[4]
port 9 nsew
flabel metal3 s -19 177 -13 183 7 FreeSans 24 0 0 0 pin_input[5]
port 10 nsew
flabel metal2 s 1549 2037 1555 2043 3 FreeSans 24 90 0 0 pin_input[6]
port 11 nsew
flabel metal2 s 1485 2037 1491 2043 3 FreeSans 24 90 0 0 pin_input[7]
port 12 nsew
flabel metal3 s 2973 977 2979 983 3 FreeSans 24 0 0 0 pin_input[8]
port 13 nsew
flabel metal2 s 781 2037 787 2043 3 FreeSans 24 90 0 0 pin_input[9]
port 14 nsew
flabel metal2 s 1245 2037 1251 2043 3 FreeSans 24 90 0 0 pin_input[10]
port 15 nsew
flabel metal3 s -19 837 -13 843 7 FreeSans 24 0 0 0 pin_input[11]
port 16 nsew
flabel metal3 s 2973 557 2979 563 3 FreeSans 24 0 0 0 pin_input[12]
port 17 nsew
flabel metal2 s 2221 2037 2227 2043 3 FreeSans 24 90 0 0 pin_input[13]
port 18 nsew
flabel metal2 s 2525 2037 2531 2043 3 FreeSans 24 90 0 0 pin_input[14]
port 19 nsew
flabel metal3 s -19 1537 -13 1543 7 FreeSans 24 0 0 0 pin_input[15]
port 20 nsew
flabel metal2 s 1085 2037 1091 2043 3 FreeSans 24 90 0 0 correct_pin
port 21 nsew
flabel metal3 s -19 1457 -13 1463 7 FreeSans 24 0 0 0 balance_check
port 22 nsew
flabel metal3 s -19 1497 -13 1503 7 FreeSans 24 0 0 0 withdraw
port 23 nsew
flabel metal3 s -19 1697 -13 1703 7 FreeSans 24 0 0 0 print_balance
port 24 nsew
flabel metal3 s -19 1897 -13 1903 7 FreeSans 24 0 0 0 amount_entered
port 25 nsew
flabel metal2 s 493 2037 499 2043 3 FreeSans 24 90 0 0 cash_eject
port 26 nsew
flabel metal3 s -19 1937 -13 1943 7 FreeSans 24 0 0 0 exit
port 27 nsew
flabel metal3 s -19 1297 -13 1303 7 FreeSans 24 0 0 0 state[0]
port 28 nsew
flabel metal2 s 381 2037 387 2043 3 FreeSans 24 90 0 0 state[1]
port 29 nsew
flabel metal2 s 653 2037 659 2043 3 FreeSans 24 90 0 0 state[2]
port 30 nsew
flabel metal2 s 1277 2037 1283 2043 3 FreeSans 24 90 0 0 auth_success
port 31 nsew
flabel metal2 s 1133 -23 1139 -17 7 FreeSans 24 270 0 0 freeze
port 32 nsew
<< end >>
