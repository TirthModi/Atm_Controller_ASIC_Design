* NGSPICE file created from atm_fsm.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR Q CLK R S D gnd vdd
.ends

* Black-box entry subcircuit for BUFX4 abstract view
.subckt BUFX4 A gnd Y vdd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A gnd Y vdd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A gnd Y vdd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C gnd Y vdd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B gnd Y vdd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D gnd Y vdd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B gnd Y vdd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A gnd Y vdd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A gnd Y vdd
.ends

.subckt atm_fsm vdd gnd clk reset insert_card pin_input[0] pin_input[1] pin_input[2]
+ pin_input[3] pin_input[4] pin_input[5] pin_input[6] pin_input[7] pin_input[8] pin_input[9]
+ pin_input[10] pin_input[11] pin_input[12] pin_input[13] pin_input[14] pin_input[15]
+ correct_pin balance_check withdraw print_balance amount_entered cash_eject exit
+ state[0] state[1] state[2] auth_success freeze
XFILL_0_0_2 gnd vdd FILL
XNOR2X1_26 BUFX4_8/Y NOR2X1_26/B gnd DFFSR_31/D vdd NOR2X1
XFILL_1_1_0 gnd vdd FILL
XBUFX2_3 BUFX2_3/A gnd auth_success vdd BUFX2
XFILL_9_1 gnd vdd FILL
XFILL_7_0_2 gnd vdd FILL
XNAND3X1_18 DFFSR_21/Q BUFX4_14/Y BUFX2_2/Y gnd NAND3X1_18/Y vdd NAND3X1
XOAI21X1_34 BUFX4_3/Y NOR2X1_3/B NOR2X1_8/A gnd NOR2X1_28/B vdd OAI21X1
XOAI22X1_1 BUFX4_7/Y OAI22X1_1/B INVX2_7/Y OR2X2_2/B gnd DFFSR_6/D vdd OAI22X1
XNAND2X1_13 INVX1_9/Y INVX1_8/Y gnd NAND2X1_14/B vdd NAND2X1
XFILL_8_1_0 gnd vdd FILL
XNAND2X1_2 INVX1_2/Y NOR2X1_2/Y gnd NOR2X1_3/B vdd NAND2X1
XNOR2X1_27 BUFX4_8/Y NOR2X1_27/B gnd DFFSR_32/D vdd NOR2X1
XDFFSR_19 DFFSR_19/Q CLKBUF1_6/Y DFFSR_5/R vdd DFFSR_19/D gnd vdd DFFSR
XFILL_1_1_1 gnd vdd FILL
XBUFX2_4 BUFX2_4/A gnd freeze vdd BUFX2
XOAI21X1_35 BUFX4_3/Y NOR2X1_3/B DFFSR_34/Q gnd NOR2X1_29/B vdd OAI21X1
XNAND2X1_14 XNOR2X1_2/A NAND2X1_14/B gnd OAI21X1_9/A vdd NAND2X1
XFILL_8_1_1 gnd vdd FILL
XFILL_9_2 gnd vdd FILL
XNAND2X1_3 DFFSR_24/Q AND2X2_2/Y gnd NAND2X1_3/Y vdd NAND2X1
XNAND3X1_19 DFFSR_22/Q BUFX4_14/Y BUFX4_1/Y gnd OAI21X1_23/C vdd NAND3X1
XOAI22X1_2 INVX1_3/Y INVX2_8/Y NOR2X1_36/Y OAI22X1_2/D gnd OAI22X1_2/Y vdd OAI22X1
XBUFX4_10 BUFX4_8/A gnd BUFX2_4/A vdd BUFX4
XNOR2X1_28 BUFX4_8/Y NOR2X1_28/B gnd DFFSR_33/D vdd NOR2X1
XDFFSR_20 INVX2_6/A CLKBUF1_4/Y DFFSR_23/R vdd DFFSR_20/D gnd vdd DFFSR
XFILL_1_1_2 gnd vdd FILL
XXOR2X1_1 XOR2X1_1/A DFFSR_10/Q gnd XOR2X1_1/Y vdd XOR2X1
XNAND3X1_20 DFFSR_22/Q DFFSR_21/Q NOR2X1_19/Y gnd NAND2X1_18/B vdd NAND3X1
XOAI21X1_36 BUFX4_3/Y NOR2X1_3/B NOR2X1_7/A gnd NOR2X1_30/B vdd OAI21X1
XNAND2X1_4 NOR2X1_7/Y NOR2X1_8/Y gnd NAND2X1_4/Y vdd NAND2X1
XNAND2X1_15 NOR3X1_2/C OAI21X1_11/Y gnd NAND2X1_15/Y vdd NAND2X1
XBUFX2_5 BUFX2_5/A gnd state[0] vdd BUFX2
XFILL_8_1_2 gnd vdd FILL
XDFFSR_21 DFFSR_21/Q CLKBUF1_6/Y DFFSR_5/R vdd DFFSR_21/D gnd vdd DFFSR
XBUFX4_11 INVX8_1/Y gnd BUFX4_11/Y vdd BUFX4
XNOR2X1_29 BUFX4_8/Y NOR2X1_29/B gnd DFFSR_34/D vdd NOR2X1
XNAND2X1_16 OAI21X1_14/Y INVX1_10/Y gnd NAND2X1_16/Y vdd NAND2X1
XFILL_4_0_0 gnd vdd FILL
XOAI21X1_37 BUFX4_5/Y NOR2X1_3/B DFFSR_36/Q gnd NOR2X1_31/B vdd OAI21X1
XINVX2_1 BUFX2_5/A gnd INVX2_1/Y vdd INVX2
XBUFX2_6 DFFSR_2/Q gnd state[1] vdd BUFX2
XNAND3X1_21 DFFSR_23/Q BUFX4_14/Y BUFX4_1/Y gnd OAI21X1_24/C vdd NAND3X1
XNAND2X1_5 NOR2X1_9/Y NOR2X1_10/Y gnd NOR2X1_11/B vdd NAND2X1
XDFFSR_22 DFFSR_22/Q CLKBUF1_6/Y DFFSR_23/R vdd DFFSR_22/D gnd vdd DFFSR
XNOR2X1_30 BUFX4_8/Y NOR2X1_30/B gnd DFFSR_35/D vdd NOR2X1
XBUFX4_12 INVX8_1/Y gnd BUFX4_12/Y vdd BUFX4
XFILL_4_0_1 gnd vdd FILL
XNAND2X1_17 NOR3X1_3/C INVX2_5/Y gnd OAI21X1_18/B vdd NAND2X1
XNAND2X1_6 NAND2X1_6/A NOR2X1_13/Y gnd NOR2X1_16/A vdd NAND2X1
XOAI21X1_38 BUFX4_6/Y NOR2X1_3/B DFFSR_37/Q gnd NOR2X1_32/B vdd OAI21X1
XINVX2_2 INVX2_2/A gnd INVX2_2/Y vdd INVX2
XBUFX2_7 INVX1_1/A gnd state[2] vdd BUFX2
XDFFSR_23 DFFSR_23/Q CLKBUF1_6/Y DFFSR_23/R vdd DFFSR_23/D gnd vdd DFFSR
XNAND3X1_22 DFFSR_21/Q AND2X2_2/Y NOR2X1_19/Y gnd NAND2X1_19/B vdd NAND3X1
XBUFX4_13 INVX8_1/Y gnd BUFX4_13/Y vdd BUFX4
XNOR2X1_31 BUFX4_9/Y NOR2X1_31/B gnd DFFSR_36/D vdd NOR2X1
XFILL_4_0_2 gnd vdd FILL
XINVX2_3 INVX2_3/A gnd INVX2_3/Y vdd INVX2
XOAI21X1_39 BUFX4_5/Y NOR2X1_3/B NOR2X1_9/B gnd NOR2X1_33/B vdd OAI21X1
XNOR2X1_1 DFFSR_2/Q INVX2_1/Y gnd NOR2X1_1/Y vdd NOR2X1
XNAND3X1_23 DFFSR_24/Q BUFX4_14/Y BUFX4_1/Y gnd OAI21X1_25/C vdd NAND3X1
XNAND2X1_18 INVX2_5/Y NAND2X1_18/B gnd NAND2X1_18/Y vdd NAND2X1
XNAND2X1_7 NOR2X1_14/Y NOR2X1_15/Y gnd NAND2X1_7/Y vdd NAND2X1
XFILL_5_1_0 gnd vdd FILL
XDFFSR_24 DFFSR_24/Q CLKBUF1_6/Y DFFSR_23/R vdd DFFSR_24/D gnd vdd DFFSR
XBUFX4_14 INVX8_1/Y gnd BUFX4_14/Y vdd BUFX4
XNOR2X1_32 BUFX4_7/Y NOR2X1_32/B gnd DFFSR_37/D vdd NOR2X1
XNAND2X1_19 INVX2_5/Y NAND2X1_19/B gnd NAND2X1_19/Y vdd NAND2X1
XOAI21X1_40 BUFX4_5/Y NOR2X1_3/B DFFSR_39/Q gnd NOR2X1_34/B vdd OAI21X1
XFILL_5_1_1 gnd vdd FILL
XNOR2X1_2 DFFSR_6/Q INVX1_3/Y gnd NOR2X1_2/Y vdd NOR2X1
XINVX2_4 INVX2_4/A gnd INVX2_4/Y vdd INVX2
XDFFSR_25 DFFSR_25/Q CLKBUF1_5/Y DFFSR_27/R vdd DFFSR_25/D gnd vdd DFFSR
XNAND2X1_8 AND2X2_3/Y NAND2X1_8/B gnd OR2X2_2/B vdd NAND2X1
XBUFX4_15 INVX8_3/Y gnd DFFSR_2/R vdd BUFX4
XNAND3X1_24 correct_pin BUFX4_11/Y INVX2_8/Y gnd AOI22X1_1/D vdd NAND3X1
XNOR2X1_33 BUFX4_7/Y NOR2X1_33/B gnd DFFSR_38/D vdd NOR2X1
XOR2X2_1 DFFSR_8/Q OR2X2_1/B gnd OR2X2_1/Y vdd OR2X2
XINVX2_5 OR2X2_2/B gnd INVX2_5/Y vdd INVX2
XOAI21X1_41 correct_pin BUFX4_6/Y INVX2_7/Y gnd OAI21X1_42/C vdd OAI21X1
XNAND2X1_9 DFFSR_8/Q OR2X2_1/B gnd XOR2X1_1/A vdd NAND2X1
XFILL_5_1_2 gnd vdd FILL
XNOR2X1_3 BUFX4_5/Y NOR2X1_3/B gnd INVX8_2/A vdd NOR2X1
XNAND3X1_25 DFFSR_2/Q INVX1_20/Y INVX1_21/Y gnd OAI21X1_52/C vdd NAND3X1
XNAND2X1_20 INVX1_2/Y INVX2_8/Y gnd OAI22X1_2/D vdd NAND2X1
XDFFSR_26 DFFSR_26/Q CLKBUF1_6/Y DFFSR_5/R vdd DFFSR_26/D gnd vdd DFFSR
XOR2X2_2 OR2X2_2/A OR2X2_2/B gnd OR2X2_2/Y vdd OR2X2
XNOR2X1_34 BUFX4_7/Y NOR2X1_34/B gnd DFFSR_39/D vdd NOR2X1
XBUFX4_16 INVX8_3/Y gnd DFFSR_7/R vdd BUFX4
XFILL_1_0_0 gnd vdd FILL
XINVX2_6 INVX2_6/A gnd INVX2_6/Y vdd INVX2
XNOR2X1_4 DFFSR_21/Q DFFSR_19/Q gnd NOR2X1_4/Y vdd NOR2X1
XOAI21X1_42 INVX2_7/Y BUFX4_6/Y OAI21X1_42/C gnd OAI22X1_1/B vdd OAI21X1
XFILL_8_1 gnd vdd FILL
XNAND2X1_21 BUFX4_11/Y OAI22X1_2/Y gnd OAI21X1_43/C vdd NAND2X1
XDFFSR_27 DFFSR_27/Q CLKBUF1_5/Y DFFSR_27/R vdd DFFSR_27/D gnd vdd DFFSR
XINVX1_10 INVX1_10/A gnd INVX1_10/Y vdd INVX1
XBUFX4_17 INVX8_3/Y gnd DFFSR_8/R vdd BUFX4
XFILL_8_0_0 gnd vdd FILL
XNOR2X1_35 INVX1_3/A INVX2_7/Y gnd NOR2X1_35/Y vdd NOR2X1
XOR2X2_3 OR2X2_3/A OR2X2_3/B gnd OR2X2_3/Y vdd OR2X2
XFILL_1_0_1 gnd vdd FILL
XINVX2_7 DFFSR_6/Q gnd INVX2_7/Y vdd INVX2
XAOI21X1_1 NOR2X1_6/Y AND2X2_1/Y NAND2X1_3/Y gnd OAI21X1_2/C vdd AOI21X1
XNOR2X1_5 INVX1_6/Y INVX2_2/Y gnd NOR2X1_6/B vdd NOR2X1
XFILL_8_2 gnd vdd FILL
XOAI21X1_43 INVX1_3/Y OR2X2_2/B OAI21X1_43/C gnd DFFSR_7/D vdd OAI21X1
XNAND2X1_22 INVX2_9/Y INVX2_1/Y gnd NOR2X1_37/B vdd NAND2X1
XFILL_8_0_1 gnd vdd FILL
XBUFX4_18 INVX8_3/Y gnd DFFSR_5/R vdd BUFX4
XINVX1_11 INVX1_11/A gnd INVX1_11/Y vdd INVX1
XDFFSR_28 DFFSR_28/Q CLKBUF1_2/Y DFFSR_2/R vdd DFFSR_28/D gnd vdd DFFSR
XNAND3X1_1 DFFSR_8/Q BUFX4_13/Y BUFX4_2/Y gnd OAI21X1_3/C vdd NAND3X1
XNOR2X1_36 NOR2X1_2/Y NOR2X1_35/Y gnd NOR2X1_36/Y vdd NOR2X1
XFILL_1_0_2 gnd vdd FILL
XFILL_2_1_0 gnd vdd FILL
XAOI21X1_2 INVX1_10/A INVX1_11/A DFFSR_19/Q gnd AOI21X1_2/Y vdd AOI21X1
XOAI21X1_44 BUFX4_7/Y BUFX2_2/Y OR2X2_2/B gnd DFFSR_5/D vdd OAI21X1
XNOR2X1_6 NOR2X1_6/A NOR2X1_6/B gnd NOR2X1_6/Y vdd NOR2X1
XFILL_8_3 gnd vdd FILL
XINVX2_8 BUFX4_6/Y gnd INVX2_8/Y vdd INVX2
XNAND2X1_23 INVX2_1/Y INVX1_16/A gnd INVX1_18/A vdd NAND2X1
XINVX1_12 DFFSR_21/Q gnd INVX1_12/Y vdd INVX1
XDFFSR_29 DFFSR_29/Q CLKBUF1_2/Y DFFSR_2/R vdd DFFSR_29/D gnd vdd DFFSR
XFILL_9_1_0 gnd vdd FILL
XFILL_8_0_2 gnd vdd FILL
XNAND3X1_2 INVX2_6/A INVX1_11/A INVX2_3/Y gnd NOR2X1_6/A vdd NAND3X1
XBUFX4_19 INVX8_3/Y gnd DFFSR_23/R vdd BUFX4
XNOR2X1_37 INVX1_1/A NOR2X1_37/B gnd NOR2X1_37/Y vdd NOR2X1
XINVX2_9 DFFSR_2/Q gnd INVX2_9/Y vdd INVX2
XAOI21X1_3 OR2X2_2/A DFFSR_22/Q DFFSR_23/Q gnd AOI21X1_3/Y vdd AOI21X1
XFILL_2_1_1 gnd vdd FILL
XNOR2X1_7 NOR2X1_7/A DFFSR_34/Q gnd NOR2X1_7/Y vdd NOR2X1
XNAND2X1_24 INVX1_17/Y NOR2X1_39/Y gnd NAND2X1_24/Y vdd NAND2X1
XINVX1_1 INVX1_1/A gnd INVX1_1/Y vdd INVX1
XOAI21X1_45 NOR2X1_2/Y OAI22X1_2/D BUFX4_11/Y gnd NOR2X1_42/A vdd OAI21X1
XINVX1_13 INVX1_13/A gnd INVX1_13/Y vdd INVX1
XDFFSR_30 DFFSR_30/Q CLKBUF1_4/Y DFFSR_5/R vdd DFFSR_30/D gnd vdd DFFSR
XBUFX4_20 INVX8_3/Y gnd DFFSR_27/R vdd BUFX4
XNAND3X1_3 OR2X2_1/B BUFX4_13/Y BUFX4_2/Y gnd NAND3X1_3/Y vdd NAND3X1
XFILL_9_1_1 gnd vdd FILL
XNOR2X1_38 INVX1_1/A INVX2_9/Y gnd INVX1_16/A vdd NOR2X1
XNOR2X1_8 NOR2X1_8/A DFFSR_32/Q gnd NOR2X1_8/Y vdd NOR2X1
XAOI21X1_4 OR2X2_2/A AND2X2_2/Y DFFSR_24/Q gnd AOI21X1_4/Y vdd AOI21X1
XOAI21X1_10 XNOR2X1_2/Y OR2X2_2/B NAND3X1_9/Y gnd DFFSR_14/D vdd OAI21X1
XOAI21X1_46 amount_entered NOR2X1_39/Y NOR2X1_40/Y gnd OAI21X1_47/C vdd OAI21X1
XNAND2X1_25 INVX1_1/A INVX2_1/Y gnd INVX1_21/A vdd NAND2X1
XFILL_2_1_2 gnd vdd FILL
XINVX1_14 BUFX2_3/A gnd INVX1_14/Y vdd INVX1
XFILL_9_1_2 gnd vdd FILL
XINVX1_2 correct_pin gnd INVX1_2/Y vdd INVX1
XDFFSR_31 DFFSR_31/Q CLKBUF1_2/Y DFFSR_2/R vdd DFFSR_31/D gnd vdd DFFSR
XNOR2X1_39 exit INVX2_1/Y gnd NOR2X1_39/Y vdd NOR2X1
XNAND3X1_4 DFFSR_10/Q BUFX4_13/Y BUFX4_2/Y gnd OAI21X1_5/C vdd NAND3X1
XFILL_3_1 gnd vdd FILL
XNOR2X1_9 DFFSR_39/Q NOR2X1_9/B gnd NOR2X1_9/Y vdd NOR2X1
XOAI21X1_11 INVX2_2/Y XNOR2X1_2/A INVX1_6/Y gnd OAI21X1_11/Y vdd OAI21X1
XINVX1_3 INVX1_3/A gnd INVX1_3/Y vdd INVX1
XAOI21X1_5 INVX2_1/Y BUFX4_9/Y AOI21X1_5/C gnd DFFSR_1/D vdd AOI21X1
XDFFSR_1 BUFX2_5/A CLKBUF1_2/Y DFFSR_2/R vdd DFFSR_1/D gnd vdd DFFSR
XNAND2X1_26 insert_card NOR2X1_37/Y gnd OAI21X1_48/C vdd NAND2X1
XOAI21X1_47 INVX1_16/Y NAND2X1_24/Y OAI21X1_47/C gnd NOR2X1_41/B vdd OAI21X1
XDFFSR_32 DFFSR_32/Q CLKBUF1_5/Y DFFSR_27/R vdd DFFSR_32/D gnd vdd DFFSR
XFILL_5_0_0 gnd vdd FILL
XINVX1_15 balance_check gnd INVX1_15/Y vdd INVX1
XNOR2X1_40 DFFSR_2/Q INVX1_21/A gnd NOR2X1_40/Y vdd NOR2X1
XNAND3X1_5 INVX2_4/A BUFX4_13/Y BUFX2_1/Y gnd NAND3X1_5/Y vdd NAND3X1
XDFFSR_2 DFFSR_2/Q CLKBUF1_2/Y DFFSR_2/R vdd DFFSR_2/D gnd vdd DFFSR
XOAI21X1_12 NAND2X1_15/Y OR2X2_2/B OAI21X1_12/C gnd DFFSR_15/D vdd OAI21X1
XOAI21X1_48 cash_eject NAND2X1_27/Y OAI21X1_48/C gnd NOR2X1_41/A vdd OAI21X1
XNAND2X1_27 INVX1_1/A NOR2X1_1/Y gnd NAND2X1_27/Y vdd NAND2X1
XINVX1_4 INVX1_4/A gnd INVX1_4/Y vdd INVX1
XFILL_5_0_1 gnd vdd FILL
XINVX1_16 INVX1_16/A gnd INVX1_16/Y vdd INVX1
XAOI21X1_6 AOI21X1_6/A INVX1_19/A BUFX4_9/Y gnd AOI22X1_3/D vdd AOI21X1
XNAND3X1_6 DFFSR_8/Q DFFSR_10/Q OR2X2_1/B gnd NOR3X1_1/C vdd NAND3X1
XDFFSR_33 NOR2X1_8/A CLKBUF1_5/Y DFFSR_27/R vdd DFFSR_33/D gnd vdd DFFSR
XNOR2X1_41 NOR2X1_41/A NOR2X1_41/B gnd NOR2X1_41/Y vdd NOR2X1
XINVX1_5 INVX1_5/A gnd INVX1_5/Y vdd INVX1
XOAI21X1_13 XNOR2X1_3/Y OR2X2_2/B OAI21X1_13/C gnd DFFSR_16/D vdd OAI21X1
XDFFSR_3 INVX1_1/A CLKBUF1_1/Y DFFSR_7/R vdd DFFSR_3/D gnd vdd DFFSR
XNAND2X1_28 BUFX2_5/A INVX1_16/A gnd NAND2X1_28/Y vdd NAND2X1
XOAI21X1_49 INVX1_15/Y INVX1_18/A NOR2X1_41/Y gnd NOR2X1_42/B vdd OAI21X1
XDFFSR_34 DFFSR_34/Q CLKBUF1_5/Y DFFSR_27/R vdd DFFSR_34/D gnd vdd DFFSR
XFILL_5_0_2 gnd vdd FILL
XFILL_6_1_0 gnd vdd FILL
XINVX1_17 print_balance gnd INVX1_17/Y vdd INVX1
XNOR3X1_1 INVX1_7/Y INVX2_4/Y NOR3X1_1/C gnd INVX1_8/A vdd NOR3X1
XNAND3X1_7 INVX1_7/A BUFX4_13/Y BUFX2_1/Y gnd OAI21X1_8/C vdd NAND3X1
XNOR2X1_42 NOR2X1_42/A NOR2X1_42/B gnd AOI21X1_5/C vdd NOR2X1
XOAI21X1_50 exit INVX2_9/Y INVX1_17/Y gnd INVX1_19/A vdd OAI21X1
XAND2X2_1 NOR2X1_4/Y INVX1_5/Y gnd AND2X2_1/Y vdd AND2X2
XOAI21X1_14 INVX2_3/Y NOR3X1_2/C INVX1_5/Y gnd OAI21X1_14/Y vdd OAI21X1
XINVX1_6 INVX1_6/A gnd INVX1_6/Y vdd INVX1
XDFFSR_4 BUFX2_3/A CLKBUF1_1/Y DFFSR_7/R vdd DFFSR_4/D gnd vdd DFFSR
XDFFSR_35 NOR2X1_7/A CLKBUF1_5/Y DFFSR_27/R vdd DFFSR_35/D gnd vdd DFFSR
XNOR3X1_2 INVX1_5/Y INVX2_3/Y NOR3X1_2/C gnd INVX1_10/A vdd NOR3X1
XFILL_6_1_1 gnd vdd FILL
XNAND3X1_8 INVX1_9/A BUFX4_13/Y BUFX2_1/Y gnd OAI21X1_9/C vdd NAND3X1
XNOR2X1_43 INVX1_18/A NOR2X1_43/B gnd NOR2X1_43/Y vdd NOR2X1
XINVX1_18 INVX1_18/A gnd INVX1_18/Y vdd INVX1
XAND2X2_2 DFFSR_23/Q DFFSR_22/Q gnd AND2X2_2/Y vdd AND2X2
XDFFSR_5 BUFX4_8/A CLKBUF1_4/Y DFFSR_5/R vdd DFFSR_5/D gnd vdd DFFSR
XOAI21X1_15 OR2X2_2/B NAND2X1_16/Y NAND3X1_13/Y gnd DFFSR_17/D vdd OAI21X1
XINVX1_7 INVX1_7/A gnd INVX1_7/Y vdd INVX1
XOAI21X1_51 withdraw INVX1_19/Y INVX1_15/Y gnd AOI22X1_2/D vdd OAI21X1
XNOR3X1_3 INVX1_12/Y INVX2_6/Y NOR3X1_3/C gnd OR2X2_2/A vdd NOR3X1
XDFFSR_36 DFFSR_36/Q CLKBUF1_2/Y DFFSR_2/R vdd DFFSR_36/D gnd vdd DFFSR
XFILL_6_1_2 gnd vdd FILL
XINVX1_19 INVX1_19/A gnd INVX1_19/Y vdd INVX1
XBUFX4_1 BUFX2_2/A gnd BUFX4_1/Y vdd BUFX4
XNAND3X1_9 INVX2_2/A BUFX4_12/Y BUFX2_1/Y gnd NAND3X1_9/Y vdd NAND3X1
XOAI21X1_52 INVX2_1/Y INVX1_16/Y OAI21X1_52/C gnd AOI21X1_6/A vdd OAI21X1
XAND2X2_3 AND2X2_3/A AND2X2_3/B gnd AND2X2_3/Y vdd AND2X2
XOAI21X1_16 INVX1_11/Y INVX1_10/Y INVX2_5/Y gnd OAI21X1_17/B vdd OAI21X1
XDFFSR_6 DFFSR_6/Q CLKBUF1_4/Y DFFSR_5/R vdd DFFSR_6/D gnd vdd DFFSR
XINVX1_8 INVX1_8/A gnd INVX1_8/Y vdd INVX1
XFILL_2_0_0 gnd vdd FILL
XDFFSR_37 DFFSR_37/Q CLKBUF1_1/Y DFFSR_7/R vdd DFFSR_37/D gnd vdd DFFSR
XINVX1_20 exit gnd INVX1_20/Y vdd INVX1
XFILL_9_0_0 gnd vdd FILL
XBUFX4_2 BUFX2_2/A gnd BUFX4_2/Y vdd BUFX4
XOAI21X1_17 NOR2X1_17/Y OAI21X1_17/B OAI21X1_17/C gnd DFFSR_18/D vdd OAI21X1
XINVX1_9 INVX1_9/A gnd INVX1_9/Y vdd INVX1
XOAI21X1_53 exit INVX1_1/Y INVX1_17/Y gnd INVX1_22/A vdd OAI21X1
XDFFSR_7 INVX1_3/A CLKBUF1_1/Y DFFSR_7/R vdd DFFSR_7/D gnd vdd DFFSR
XFILL_2_0_1 gnd vdd FILL
XAND2X2_4 NOR3X1_3/C INVX2_6/Y gnd AND2X2_4/Y vdd AND2X2
XDFFSR_38 NOR2X1_9/B CLKBUF1_1/Y DFFSR_7/R vdd DFFSR_38/D gnd vdd DFFSR
XINVX1_21 INVX1_21/A gnd INVX1_21/Y vdd INVX1
XAOI22X1_1 BUFX4_11/Y NOR2X1_37/Y INVX1_14/Y AOI22X1_1/D gnd DFFSR_4/D vdd AOI22X1
XBUFX4_3 BUFX4_3/A gnd BUFX4_3/Y vdd BUFX4
XNOR2X1_10 DFFSR_37/Q DFFSR_36/Q gnd NOR2X1_10/Y vdd NOR2X1
XFILL_9_0_1 gnd vdd FILL
XXNOR2X1_1 NOR3X1_1/C INVX2_4/Y gnd OAI21X1_6/A vdd XNOR2X1
XOAI21X1_18 AOI21X1_2/Y OAI21X1_18/B NAND3X1_15/Y gnd DFFSR_19/D vdd OAI21X1
XDFFSR_8 DFFSR_8/Q CLKBUF1_3/Y DFFSR_8/R vdd DFFSR_8/D gnd vdd DFFSR
XOAI21X1_54 withdraw INVX1_22/A INVX1_15/Y gnd NOR2X1_43/B vdd OAI21X1
XFILL_2_0_2 gnd vdd FILL
XFILL_3_1_0 gnd vdd FILL
XDFFSR_39 DFFSR_39/Q CLKBUF1_2/Y DFFSR_2/R vdd DFFSR_39/D gnd vdd DFFSR
XFILL_9_0_2 gnd vdd FILL
XINVX1_22 INVX1_22/A gnd INVX1_22/Y vdd INVX1
XAOI22X1_2 correct_pin INVX2_8/Y INVX1_18/Y AOI22X1_2/D gnd AOI22X1_3/C vdd AOI22X1
XNOR2X1_11 NAND2X1_4/Y NOR2X1_11/B gnd AND2X2_3/B vdd NOR2X1
XBUFX4_4 BUFX4_3/A gnd BUFX4_4/Y vdd BUFX4
XXNOR2X1_2 XNOR2X1_2/A INVX2_2/Y gnd XNOR2X1_2/Y vdd XNOR2X1
XOAI21X1_19 INVX2_6/Y NOR3X1_3/C INVX2_5/Y gnd OAI21X1_19/Y vdd OAI21X1
XOAI21X1_55 INVX1_20/Y amount_entered NOR2X1_40/Y gnd OAI21X1_56/C vdd OAI21X1
XDFFSR_9 OR2X2_1/B CLKBUF1_3/Y DFFSR_8/R vdd DFFSR_9/D gnd vdd DFFSR
XFILL_3_1_1 gnd vdd FILL
XNOR2X1_12 DFFSR_31/Q DFFSR_30/Q gnd NAND2X1_6/A vdd NOR2X1
XBUFX4_5 BUFX4_3/A gnd BUFX4_5/Y vdd BUFX4
XXNOR2X1_3 NOR3X1_2/C INVX2_3/Y gnd XNOR2X1_3/Y vdd XNOR2X1
XAOI22X1_3 INVX2_9/Y BUFX4_9/Y AOI22X1_3/C AOI22X1_3/D gnd DFFSR_2/D vdd AOI22X1
XOAI21X1_20 AND2X2_4/Y OAI21X1_19/Y OAI21X1_20/C gnd DFFSR_20/D vdd OAI21X1
XOAI21X1_56 NAND2X1_28/Y INVX1_22/Y OAI21X1_56/C gnd OR2X2_3/A vdd OAI21X1
XFILL_3_1_2 gnd vdd FILL
XNOR2X1_13 DFFSR_29/Q DFFSR_28/Q gnd NOR2X1_13/Y vdd NOR2X1
XBUFX4_6 BUFX4_3/A gnd BUFX4_6/Y vdd BUFX4
XOAI21X1_21 INVX2_6/Y NOR3X1_3/C INVX1_12/Y gnd INVX1_13/A vdd OAI21X1
XOAI21X1_57 cash_eject NAND2X1_27/Y OAI21X1_52/C gnd OR2X2_3/B vdd OAI21X1
XNOR2X1_14 DFFSR_27/Q DFFSR_26/Q gnd NOR2X1_14/Y vdd NOR2X1
XFILL_6_0_0 gnd vdd FILL
XBUFX4_7 BUFX4_8/A gnd BUFX4_7/Y vdd BUFX4
XOAI21X1_22 INVX1_13/Y OR2X2_2/Y NAND3X1_18/Y gnd DFFSR_21/D vdd OAI21X1
XOAI21X1_58 NOR2X1_43/Y OR2X2_3/Y BUFX4_11/Y gnd OAI21X1_58/Y vdd OAI21X1
XFILL_6_1 gnd vdd FILL
XCLKBUF1_1 clk gnd CLKBUF1_1/Y vdd CLKBUF1
XNOR2X1_15 DFFSR_25/Q BUFX4_14/Y gnd NOR2X1_15/Y vdd NOR2X1
XBUFX4_8 BUFX4_8/A gnd BUFX4_8/Y vdd BUFX4
XFILL_6_0_1 gnd vdd FILL
XOAI21X1_59 INVX1_1/Y BUFX4_11/Y OAI21X1_58/Y gnd DFFSR_3/D vdd OAI21X1
XOAI21X1_23 NOR2X1_18/Y NAND2X1_18/Y OAI21X1_23/C gnd DFFSR_22/D vdd OAI21X1
XCLKBUF1_2 clk gnd CLKBUF1_2/Y vdd CLKBUF1
XFILL_0_1_0 gnd vdd FILL
XNOR2X1_16 NOR2X1_16/A NAND2X1_7/Y gnd AND2X2_3/A vdd NOR2X1
XFILL_6_2 gnd vdd FILL
XFILL_6_0_2 gnd vdd FILL
XBUFX4_9 BUFX4_8/A gnd BUFX4_9/Y vdd BUFX4
XFILL_7_1_0 gnd vdd FILL
XOAI21X1_24 AOI21X1_3/Y NAND2X1_19/Y OAI21X1_24/C gnd DFFSR_23/D vdd OAI21X1
XOAI21X1_1 DFFSR_19/Q INVX1_11/A INVX2_6/A gnd INVX1_4/A vdd OAI21X1
XINVX8_1 BUFX4_7/Y gnd INVX8_1/Y vdd INVX8
XCLKBUF1_3 clk gnd CLKBUF1_3/Y vdd CLKBUF1
XFILL_0_1_1 gnd vdd FILL
XNOR2X1_17 INVX1_11/A INVX1_10/A gnd NOR2X1_17/Y vdd NOR2X1
XFILL_7_1_1 gnd vdd FILL
XFILL_10_1 gnd vdd FILL
XOAI21X1_2 DFFSR_21/Q INVX1_4/Y OAI21X1_2/C gnd NAND2X1_8/B vdd OAI21X1
XINVX8_2 INVX8_2/A gnd BUFX2_2/A vdd INVX8
XOAI21X1_25 OR2X2_2/B AOI21X1_4/Y OAI21X1_25/C gnd DFFSR_24/D vdd OAI21X1
XCLKBUF1_4 clk gnd CLKBUF1_4/Y vdd CLKBUF1
XFILL_0_1_2 gnd vdd FILL
XNOR2X1_18 DFFSR_22/Q OR2X2_2/A gnd NOR2X1_18/Y vdd NOR2X1
XDFFSR_10 DFFSR_10/Q CLKBUF1_3/Y DFFSR_8/R vdd DFFSR_10/D gnd vdd DFFSR
XFILL_7_1_2 gnd vdd FILL
XFILL_10_2 gnd vdd FILL
XOAI21X1_3 DFFSR_8/Q OR2X2_2/B OAI21X1_3/C gnd DFFSR_8/D vdd OAI21X1
XINVX8_3 reset gnd INVX8_3/Y vdd INVX8
XOAI21X1_26 BUFX4_4/Y NOR2X1_3/B DFFSR_25/Q gnd NOR2X1_20/B vdd OAI21X1
XCLKBUF1_5 clk gnd CLKBUF1_5/Y vdd CLKBUF1
XNAND3X1_10 INVX1_6/A BUFX4_12/Y BUFX4_2/Y gnd OAI21X1_12/C vdd NAND3X1
XNOR2X1_19 INVX2_6/Y NOR3X1_3/C gnd NOR2X1_19/Y vdd NOR2X1
XFILL_3_0_0 gnd vdd FILL
XDFFSR_11 INVX2_4/A CLKBUF1_3/Y DFFSR_8/R vdd DFFSR_11/D gnd vdd DFFSR
XOAI21X1_4 OAI21X1_4/A OR2X2_2/B NAND3X1_3/Y gnd DFFSR_9/D vdd OAI21X1
XCLKBUF1_6 clk gnd CLKBUF1_6/Y vdd CLKBUF1
XOAI21X1_27 BUFX4_4/Y NOR2X1_3/B DFFSR_26/Q gnd NOR2X1_21/B vdd OAI21X1
XFILL_1_1 gnd vdd FILL
XNAND3X1_11 INVX1_9/A NOR2X1_6/B INVX1_8/A gnd NOR3X1_2/C vdd NAND3X1
XDFFSR_12 INVX1_7/A CLKBUF1_1/Y DFFSR_7/R vdd DFFSR_12/D gnd vdd DFFSR
XNOR2X1_20 BUFX2_4/A NOR2X1_20/B gnd DFFSR_25/D vdd NOR2X1
XFILL_3_0_1 gnd vdd FILL
XOAI21X1_28 BUFX4_4/Y NOR2X1_3/B DFFSR_27/Q gnd NOR2X1_22/B vdd OAI21X1
XOAI21X1_5 XOR2X1_1/Y OR2X2_2/B OAI21X1_5/C gnd DFFSR_10/D vdd OAI21X1
XNAND3X1_12 INVX2_3/A BUFX4_12/Y BUFX4_2/Y gnd OAI21X1_13/C vdd NAND3X1
XNOR2X1_21 BUFX2_4/A NOR2X1_21/B gnd DFFSR_26/D vdd NOR2X1
XFILL_3_0_2 gnd vdd FILL
XDFFSR_13 INVX1_9/A CLKBUF1_3/Y DFFSR_8/R vdd DFFSR_13/D gnd vdd DFFSR
XFILL_4_1_0 gnd vdd FILL
XOAI21X1_6 OAI21X1_6/A OR2X2_2/B NAND3X1_5/Y gnd DFFSR_11/D vdd OAI21X1
XOAI21X1_29 BUFX4_5/Y NOR2X1_3/B DFFSR_28/Q gnd NOR2X1_23/B vdd OAI21X1
XNAND3X1_13 INVX1_5/A BUFX4_12/Y BUFX4_1/Y gnd NAND3X1_13/Y vdd NAND3X1
XDFFSR_14 INVX2_2/A CLKBUF1_3/Y DFFSR_8/R vdd DFFSR_14/D gnd vdd DFFSR
XNOR2X1_22 BUFX2_4/A NOR2X1_22/B gnd DFFSR_27/D vdd NOR2X1
XFILL_4_1_1 gnd vdd FILL
XOAI21X1_30 BUFX4_4/Y NOR2X1_3/B DFFSR_29/Q gnd NOR2X1_24/B vdd OAI21X1
XOAI21X1_7 INVX2_4/Y NOR3X1_1/C INVX1_7/Y gnd OAI21X1_7/Y vdd OAI21X1
XNAND3X1_14 INVX1_11/A BUFX4_12/Y BUFX2_2/Y gnd OAI21X1_17/C vdd NAND3X1
XFILL_5_1 gnd vdd FILL
XNOR2X1_23 BUFX4_9/Y NOR2X1_23/B gnd DFFSR_28/D vdd NOR2X1
XDFFSR_15 INVX1_6/A CLKBUF1_3/Y DFFSR_8/R vdd DFFSR_15/D gnd vdd DFFSR
XFILL_4_1_2 gnd vdd FILL
XOAI21X1_8 OAI21X1_8/A OR2X2_2/B OAI21X1_8/C gnd DFFSR_12/D vdd OAI21X1
XOAI21X1_31 BUFX4_4/Y NOR2X1_3/B DFFSR_30/Q gnd NOR2X1_25/B vdd OAI21X1
XNAND2X1_10 XOR2X1_1/A OR2X2_1/Y gnd OAI21X1_4/A vdd NAND2X1
XNAND3X1_15 DFFSR_19/Q BUFX4_14/Y BUFX2_2/Y gnd NAND3X1_15/Y vdd NAND3X1
XDFFSR_16 INVX2_3/A CLKBUF1_4/Y DFFSR_23/R vdd DFFSR_16/D gnd vdd DFFSR
XFILL_0_0_0 gnd vdd FILL
XNOR2X1_24 BUFX4_8/Y NOR2X1_24/B gnd DFFSR_29/D vdd NOR2X1
XOAI21X1_32 BUFX4_3/Y NOR2X1_3/B DFFSR_31/Q gnd NOR2X1_26/B vdd OAI21X1
XBUFX2_1 BUFX2_2/A gnd BUFX2_1/Y vdd BUFX2
XOAI21X1_9 OAI21X1_9/A OR2X2_2/B OAI21X1_9/C gnd DFFSR_13/D vdd OAI21X1
XFILL_7_0_0 gnd vdd FILL
XNAND3X1_16 DFFSR_19/Q INVX1_11/A INVX1_10/A gnd NOR3X1_3/C vdd NAND3X1
XNAND2X1_11 OAI21X1_7/Y INVX1_8/Y gnd OAI21X1_8/A vdd NAND2X1
XNOR2X1_25 BUFX2_4/A NOR2X1_25/B gnd DFFSR_30/D vdd NOR2X1
XDFFSR_17 INVX1_5/A CLKBUF1_4/Y DFFSR_23/R vdd DFFSR_17/D gnd vdd DFFSR
XFILL_0_0_1 gnd vdd FILL
XOAI21X1_33 BUFX4_3/Y NOR2X1_3/B DFFSR_32/Q gnd NOR2X1_27/B vdd OAI21X1
XBUFX2_2 BUFX2_2/A gnd BUFX2_2/Y vdd BUFX2
XNAND2X1_12 INVX1_9/A INVX1_8/A gnd XNOR2X1_2/A vdd NAND2X1
XFILL_7_0_1 gnd vdd FILL
XNAND3X1_17 INVX2_6/A BUFX4_12/Y BUFX4_1/Y gnd OAI21X1_20/C vdd NAND3X1
XDFFSR_18 INVX1_11/A CLKBUF1_1/Y DFFSR_7/R vdd DFFSR_18/D gnd vdd DFFSR
XNAND2X1_1 INVX1_1/Y NOR2X1_1/Y gnd BUFX4_3/A vdd NAND2X1
.ends

